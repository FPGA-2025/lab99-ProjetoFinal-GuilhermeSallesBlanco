// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.14.0.75.2
// Netlist written on Wed Oct 08 19:45:10 2025
//
// Verilog Description of module top
//

module top (fastclk, rstn, sda, scl, led) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(5[8:11])
    input fastclk;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(6[16:23])
    input rstn;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(7[16:20])
    inout sda /* synthesis black_box_pad_pin=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(8[16:19])
    inout scl /* synthesis black_box_pad_pin=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(9[16:19])
    output [3:0]led;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(10[20:23])
    
    wire fastclk_c /* synthesis SET_AS_NETWORK=fastclk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(6[16:23])
    
    wire GND_net, VCC_net, rstn_c, led_c_3, led_c_2, led_c_1, led_c_0;
    wire [15:0]por;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(15[16:19])
    
    wire sda_t, scl_t, sda_in;
    wire [15:0]cnt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(33[16:19])
    
    wire n2741, n2740;
    wire [3:0]bitidx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(35[15:21])
    wire [7:0]tx_byte;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(36[15:22])
    wire [7:0]rx_byte;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(37[15:22])
    
    wire rx_ready;
    wire [31:0]gap;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(40[16:19])
    wire [1:0]desired_read_len;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(43[15:31])
    wire [1:0]rx_remaining;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(44[15:27])
    wire [1:0]rx_byte_idx;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(45[15:26])
    
    wire send_data_after_reg;
    wire [7:0]write_data;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(69[15:25])
    wire [7:0]reg_target;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(70[15:25])
    
    wire n28124;
    wire [7:0]msb;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(72[15:18])
    wire [7:0]lsb;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(72[20:23])
    wire [15:0]distance;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(73[16:24])
    
    wire rst_N_5, n2895, n2, n1876, fastclk_c_enable_91, n447, n449, 
        n452, n453, n3572, n486, n487, n488, n1, fastclk_c_enable_2, 
        n83, n82, n81, n80, n79, n78, n77, n76, n75, n74, 
        n73, n72, n71, n70, n69, n68, n67, n66, n65, n64, 
        n63, n62, n61, n60, n59, n58, n36664, n132, n57, rx_ready_N_322, 
        n85, n84, n83_adj_2202, n82_adj_2203, n81_adj_2204, n80_adj_2205, 
        n79_adj_2206, n78_adj_2207, n77_adj_2208, n76_adj_2209, n75_adj_2210, 
        n74_adj_2211, n73_adj_2212, n72_adj_2213, fastclk_c_enable_10, 
        n71_adj_2214, n70_adj_2215, n13, n33441, n14113, n66_adj_2216, 
        n72_adj_2217, n63_adj_2218, n90, n51, n138, n75_adj_2219, 
        n78_adj_2220, n81_adj_2221, n2748, n48, n13806, n141, n45, 
        n34268;
    wire [3:0]bitidx_3__N_195;
    wire [1:0]rx_remaining_1__N_292;
    wire [15:0]cnt_15__N_167;
    
    wire n114, n2651, n69_adj_2222, n135, n54, n3368, n36, n39, 
        n2744, n2743;
    wire [7:0]reg_target_7__N_247;
    
    wire fastclk_c_enable_36, n42, sda_t_N_296, scl_t_N_310, n111, 
        n108, n105, n102, n63_adj_2223, n126, n78_adj_2224, n99, 
        n5, n13788, n13805, n136, n75_adj_2225, n129, n60_adj_2226, 
        n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, 
        n1967, n1968, n1969, n72_adj_2227, n117, n10583, fastclk_c_enable_37, 
        fastclk_c_enable_5, n87, n96, n13803, n69_adj_2228, n120, 
        n84_adj_2229, n30511, n30510, n30509, n30570, n30508, n30507, 
        n30569, n30506, n30505, n30504, n30503, n30502, n33458, 
        n2355, n2354, n2353, n2352, n2350, n2349, n30568, n3638, 
        n66_adj_2230, n123, n30501, n66_adj_2231, fastclk_c_enable_79, 
        n81_adj_2232, n2797, n2798, n2799, n2800, n2801, n2802, 
        n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, 
        n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, 
        n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, 
        n2827, n2828, n93, n2960, fastclk_c_enable_31, fastclk_c_enable_45, 
        n30500, n3070, n3068, n30567, n30566, n13780, n68_adj_2233, 
        n71_adj_2234, n74_adj_2235, n77_adj_2236, n80_adj_2237, n83_adj_2238, 
        n86, n30499, n89, n30498, n92, n30497, n95, n30565, 
        n98, n30496, n101, n30495, n104, n30564, n107, n30493, 
        n110, n30563, n113, n30562, n116, n30480, n119, n30561, 
        n122, n125, n128, n131, n134, n137, n140, n143, n146, 
        n149, n152, n155, n158, n161, fastclk_c_enable_83, n3, 
        n39_adj_2239, n42_adj_2240, n45_adj_2241, n48_adj_2242, n51_adj_2243, 
        n54_adj_2244, n57_adj_2245, n60_adj_2246, n63_adj_2247, n66_adj_2248, 
        n69_adj_2249, n72_adj_2250, n75_adj_2251, n78_adj_2252, n81_adj_2253, 
        fastclk_c_enable_34, n33454, n38419, n58_adj_2254, fastclk_c_enable_16, 
        n45_adj_2255, n34, fastclk_c_enable_32, n33483, n34415, n30490, 
        n30488, n30486, n30485, n30483, n30477, n30481, n33398, 
        n30560, n5_adj_2256, n3_adj_2257, n56, n33457, n30559, n26, 
        n30558, n30557, n23, n20, n30479, n30478, n30494, n30556, 
        n30491, n30482, fastclk_c_enable_85, n30555, n7, n5_adj_2258, 
        n30489, n32862, n30554, n30553, n30552, n30551, n30550, 
        n38121, n33384, n30484, n30487, n30475, n30474, n30492, 
        n30473, n30472, n27974, n30471, n30549, n30548, n30470, 
        n30469, n3556, n6, n6_adj_2259, n13833, n36676, n39283, 
        fastclk_c_enable_33, n13802, n33464, n34303, n34042, fastclk_c_enable_82, 
        n38123, n38122, n38120, n38119, n36620, n38118, n38117, 
        n38116, n36614, n10614, n36610, n10610, n36608, n10608, 
        n36600, n10600, n10598, n36596, n10592, n34248, n36696, 
        n10588, n10582, n10580, n36576, n36574, n30468, fastclk_c_enable_35, 
        n36550, n36546, n36540, n36538, n36536, n36530, n36528, 
        n36522, n7_adj_2260, n36498, n36492, n13808, n36480, n36474, 
        n103, n36456, n33370, n38422, n15, n27, n36448, n36438, 
        n33465, n36428, n36426, fastclk_c_enable_15, n36422, n36418, 
        n36412, n36410, n55, n29267, n36406, n29256, n81_adj_2261, 
        n36392, n36390, n36370, n36368, n36366, n36362, n38428, 
        n33453, n34354, n38430, n33439, n33444, n33443, n30467, 
        n33442, n33440, n38429, n38427, n36684, n31205, n31204, 
        n31203, n31202, n31201, n31200, fastclk_c_enable_9, n31199, 
        n31198, n31197, n31196, n31195, n31194, n31193, n31192, 
        n38426, n38425, n30466, n33437, n38423, n34245, n27539, 
        n38421, n34410, n36672, n33469, n37787, n38420, fastclk_c_enable_14, 
        n33438, n33468, n34627, n37741, n37740, n37739, n34606, 
        n38406, n38405, n38404, n38403, n38402, n38401, n38360, 
        n38359, n38358, n38351, n38350, n38349, n38348, n38347, 
        n38346, n38345, n38344, n38343, n38342, n38341, n38340, 
        n30476, n28, n38339, n30, n38338, n38337, n38336, n38330, 
        n38329, n38328, n38327, n38326, n38325, n38324, n38323, 
        fastclk_c_enable_3, n34583, n26314, n38318, fastclk_c_enable_47, 
        n38313, n38312, n38311, n38310, n38309, n38308, n38304, 
        n34576, n38302, n38299, n34062;
    
    VHI i2 (.Z(VCC_net));
    LUT4 i1_4_lut (.A(tx_byte[7]), .B(tx_byte[6]), .C(reg_target[7]), 
         .D(reg_target[6]), .Z(n36474)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 tx_byte_7__I_0_307_i3_2_lut (.A(tx_byte[2]), .B(reg_target[2]), 
         .Z(n3_adj_2257)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam tx_byte_7__I_0_307_i3_2_lut.init = 16'h6666;
    CCU2C add_26226_4 (.A0(gap[3]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30548), 
          .COUT(n30549));
    defparam add_26226_4.INIT0 = 16'haaa0;
    defparam add_26226_4.INIT1 = 16'haaa0;
    defparam add_26226_4.INJECT1_0 = "NO";
    defparam add_26226_4.INJECT1_1 = "NO";
    CCU2C add_26226_2 (.A0(gap[0]), .B0(gap[1]), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .COUT(n30548));
    defparam add_26226_2.INIT0 = 16'h000e;
    defparam add_26226_2.INIT1 = 16'h555f;
    defparam add_26226_2.INJECT1_0 = "NO";
    defparam add_26226_2.INJECT1_1 = "NO";
    CCU2C _add_1_1298_add_4_7 (.A0(distance[6]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[7]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30492), .COUT(n30493), .S0(n66_adj_2248), 
          .S1(n63_adj_2247));
    defparam _add_1_1298_add_4_7.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_7.INJECT1_1 = "NO";
    LUT4 tx_byte_7__I_0_307_i5_2_lut (.A(tx_byte[4]), .B(reg_target[4]), 
         .Z(n5_adj_2256)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam tx_byte_7__I_0_307_i5_2_lut.init = 16'h6666;
    FD1P3IX desired_read_len_i1 (.D(n38351), .SP(fastclk_c_enable_3), .CD(n14113), 
            .CK(fastclk_c), .Q(desired_read_len[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam desired_read_len_i1.GSR = "DISABLED";
    FD1P3AX send_data_after_reg_275 (.D(n3638), .SP(fastclk_c_enable_2), 
            .CK(fastclk_c), .Q(send_data_after_reg));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam send_data_after_reg_275.GSR = "DISABLED";
    FD1S3IX rx_ready_273 (.D(rx_ready_N_322), .CK(fastclk_c), .CD(n33464), 
            .Q(rx_ready));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_ready_273.GSR = "DISABLED";
    FD1P3JX desired_read_len_i0 (.D(n38345), .SP(fastclk_c_enable_3), .PD(n14113), 
            .CK(fastclk_c), .Q(desired_read_len[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam desired_read_len_i0.GSR = "DISABLED";
    FD1P3AX rx_byte_idx__i0 (.D(n33458), .SP(fastclk_c_enable_15), .CK(fastclk_c), 
            .Q(rx_byte_idx[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte_idx__i0.GSR = "DISABLED";
    FD1P3IX rx_byte__i0 (.D(n33444), .SP(fastclk_c_enable_5), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i0.GSR = "DISABLED";
    FD1P3IX rx_remaining__i0 (.D(rx_remaining_1__N_292[0]), .SP(fastclk_c_enable_15), 
            .CD(n38323), .CK(fastclk_c), .Q(rx_remaining[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_remaining__i0.GSR = "DISABLED";
    LUT4 tx_byte_7__I_0_307_i1_2_lut (.A(tx_byte[0]), .B(reg_target[0]), 
         .Z(n1)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam tx_byte_7__I_0_307_i1_2_lut.init = 16'h6666;
    BB sda_iob (.I(GND_net), .T(sda_t), .B(sda), .O(sda_in)) /* synthesis syn_instantiated=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(24[8:58])
    CCU2C _add_1_1298_add_4_5 (.A0(distance[4]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[5]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30491), .COUT(n30492), .S0(n72_adj_2250), 
          .S1(n69_adj_2249));
    defparam _add_1_1298_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1298_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1298_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_5.INJECT1_1 = "NO";
    FD1P3IX msb__i0 (.D(rx_byte[0]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i0.GSR = "DISABLED";
    CCU2C _add_1_1298_add_4_3 (.A0(distance[2]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[3]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30490), .COUT(n30491), .S0(n78_adj_2252), 
          .S1(n75_adj_2251));
    defparam _add_1_1298_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_3.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_3.INJECT1_1 = "NO";
    FD1S3IX cnt__i0 (.D(cnt_15__N_167[0]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[0])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i0.GSR = "DISABLED";
    FD1P3IX tx_byte_i0 (.D(n2741), .SP(fastclk_c_enable_82), .CD(n38323), 
            .CK(fastclk_c), .Q(tx_byte[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i0.GSR = "DISABLED";
    FD1P3AX sda_t_268 (.D(sda_t_N_296), .SP(fastclk_c_enable_9), .CK(fastclk_c), 
            .Q(sda_t));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam sda_t_268.GSR = "DISABLED";
    BB scl_iob (.I(GND_net), .T(scl_t), .B(scl)) /* synthesis syn_instantiated=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(25[8:58])
    FD1P3AX scl_t_269 (.D(scl_t_N_310), .SP(fastclk_c_enable_10), .CK(fastclk_c), 
            .Q(scl_t));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam scl_t_269.GSR = "DISABLED";
    FD1S3IX reg_target_i0 (.D(reg_target_7__N_247[0]), .CK(fastclk_c), .CD(n38323), 
            .Q(reg_target[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i0.GSR = "DISABLED";
    FD1P3IX gap__i0 (.D(n2797), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i0.GSR = "DISABLED";
    FD1S3JX bitidx_i0 (.D(bitidx_3__N_195[0]), .CK(fastclk_c), .PD(n38323), 
            .Q(bitidx[0])) /* synthesis lse_init_val=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam bitidx_i0.GSR = "DISABLED";
    FD1S3JX bitidx_i1 (.D(bitidx_3__N_195[1]), .CK(fastclk_c), .PD(n38323), 
            .Q(bitidx[1])) /* synthesis lse_init_val=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam bitidx_i1.GSR = "DISABLED";
    FD1S3JX bitidx_i2 (.D(bitidx_3__N_195[2]), .CK(fastclk_c), .PD(n38323), 
            .Q(bitidx[2])) /* synthesis lse_init_val=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam bitidx_i2.GSR = "DISABLED";
    FD1S3IX bitidx_i3 (.D(bitidx_3__N_195[3]), .CK(fastclk_c), .CD(n38323), 
            .Q(bitidx[3])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam bitidx_i3.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_430 (.A(n36368), .B(n36370), .C(n36362), .D(n36366), 
         .Z(n15)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_430.init = 16'hfffe;
    LUT4 i1_2_lut (.A(cnt[8]), .B(cnt[10]), .Z(n36368)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3JX state_FSM_i1 (.D(n10580), .CK(fastclk_c), .PD(n38323), .Q(n1969));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i1.GSR = "DISABLED";
    FD1P3IX lsb__i0 (.D(rx_byte[0]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i0.GSR = "DISABLED";
    CCU2C _add_1_1298_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(distance[1]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30490), .S1(n81_adj_2253));
    defparam _add_1_1298_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1298_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(cnt[12]), .B(cnt[7]), .C(cnt[13]), .Z(n36370)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_adj_431 (.A(cnt[15]), .B(cnt[14]), .Z(n36362)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_431.init = 16'heeee;
    CCU2C _add_1_1292_add_4_33 (.A0(gap[31]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30489), .S0(n68_adj_2233));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_33.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_33.INIT1 = 16'h0000;
    defparam _add_1_1292_add_4_33.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_33.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_432 (.A(cnt[11]), .B(cnt[9]), .Z(n36366)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_432.init = 16'heeee;
    LUT4 i1_4_lut_adj_433 (.A(n36684), .B(tx_byte[4]), .C(n36438), .D(tx_byte[7]), 
         .Z(n33384)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut_adj_433.init = 16'hfff7;
    FD1S3JX seq_state_FSM_i1 (.D(n2349), .CK(fastclk_c), .PD(n38323), 
            .Q(n2355));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam seq_state_FSM_i1.GSR = "DISABLED";
    LUT4 i31850_2_lut (.A(tx_byte[1]), .B(tx_byte[6]), .Z(n36684)) /* synthesis lut_function=(A (B)) */ ;
    defparam i31850_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_434 (.A(tx_byte[3]), .B(tx_byte[2]), .Z(n36438)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_434.init = 16'heeee;
    CCU2C _add_1_1292_add_4_31 (.A0(gap[29]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[30]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30488), .COUT(n30489), .S0(n74_adj_2235), .S1(n71_adj_2234));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_31.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_31.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_31.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_31.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_29 (.A0(gap[27]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[28]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30487), .COUT(n30488), .S0(n80_adj_2237), .S1(n77_adj_2236));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_29.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_29.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(gap[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30474), .S1(n161));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1292_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1292_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_15 (.A0(gap[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30480), .COUT(n30481), .S0(n122), .S1(n119));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1284_add_4_17 (.A0(cnt[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30473), .S0(n36));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1284_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_13 (.A0(gap[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30479), .COUT(n30480), .S0(n128), .S1(n125));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut (.A(n1960), .B(n38312), .C(n81_adj_2261), .D(n38338), 
         .Z(fastclk_c_enable_85)) /* synthesis lut_function=(A (B+!(D))+!A !(C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_4_lut.init = 16'h8dff;
    CCU2C _add_1_1292_add_4_11 (.A0(gap[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30478), .COUT(n30479), .S0(n134), .S1(n131));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_11.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_9 (.A0(gap[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30477), .COUT(n30478), .S0(n140), .S1(n137));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_9.INJECT1_1 = "NO";
    FD1P3IX distance__i0 (.D(lsb[0]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i0.GSR = "DISABLED";
    CCU2C _add_1_1292_add_4_7 (.A0(gap[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30476), .COUT(n30477), .S0(n146), .S1(n143));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_7.INJECT1_1 = "NO";
    FD1P3AX write_data__i1 (.D(n38338), .SP(fastclk_c_enable_14), .CK(fastclk_c), 
            .Q(write_data[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam write_data__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_435 (.A(rx_byte_idx[0]), .B(n38325), .C(rx_remaining[1]), 
         .D(n38327), .Z(n33458)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_adj_435.init = 16'h8848;
    FD1P3AX por_1137__i0 (.D(n85), .SP(rst_N_5), .CK(fastclk_c), .Q(por[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i0.GSR = "DISABLED";
    CCU2C _add_1_1292_add_4_5 (.A0(gap[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30475), .COUT(n30476), .S0(n152), .S1(n149));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_3 (.A0(gap[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30474), .COUT(n30475), .S0(n158), .S1(n155));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_3.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_17 (.A0(gap[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30481), .COUT(n30482), .S0(n116), .S1(n113));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_17.INJECT1_1 = "NO";
    CCU2C _add_1_1284_add_4_15 (.A0(cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30472), .COUT(n30473), .S0(n42), .S1(n39));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_19 (.A0(gap[17]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[18]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30482), .COUT(n30483), .S0(n110), .S1(n107));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1284_add_4_13 (.A0(cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30471), .COUT(n30472), .S0(n48), .S1(n45));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n38340), .B(n38327), .C(bitidx[1]), 
         .D(bitidx[0]), .Z(n33483)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(250[21] 260[24])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_4_lut_adj_436 (.A(cnt[1]), .B(n38337), .C(cnt[6]), .D(cnt[0]), 
         .Z(n34354)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut_adj_436.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut (.A(n38327), .B(rx_remaining[1]), .C(n1960), .Z(n7)) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(271[25:38])
    defparam i1_2_lut_3_lut.init = 16'hb0b0;
    LUT4 i1_2_lut_rep_304_3_lut (.A(n38327), .B(rx_remaining[1]), .C(n1960), 
         .Z(n38309)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(271[25:38])
    defparam i1_2_lut_rep_304_3_lut.init = 16'h4040;
    LUT4 i1_3_lut_3_lut (.A(n38327), .B(n1960), .C(rx_remaining[1]), .Z(n34627)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(271[25:38])
    defparam i1_3_lut_3_lut.init = 16'h0404;
    LUT4 i1_4_lut_4_lut_adj_437 (.A(n38327), .B(n36418), .C(n37787), .D(n36498), 
         .Z(n34303)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(271[25:38])
    defparam i1_4_lut_4_lut_adj_437.init = 16'hfdfc;
    LUT4 i22363_3_lut_3_lut (.A(n38327), .B(rx_remaining[1]), .C(rx_remaining[0]), 
         .Z(n26314)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(271[25:38])
    defparam i22363_3_lut_3_lut.init = 16'hb4b4;
    GSR GSR_INST (.GSR(n38338));
    LUT4 n1837_bdd_2_lut_32394_4_lut (.A(n38327), .B(n2651), .C(n38347), 
         .D(n1965), .Z(n37787)) /* synthesis lut_function=(!(A+!(B (D)+!B !(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(271[25:38])
    defparam n1837_bdd_2_lut_32394_4_lut.init = 16'h4500;
    LUT4 i760_3_lut_4_lut (.A(n38327), .B(n38324), .C(n1964), .D(n1965), 
         .Z(n2740)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i760_3_lut_4_lut.init = 16'h3530;
    LUT4 i32185_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n27974), 
         .Z(fastclk_c_enable_37)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32185_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i32189_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n13808), 
         .Z(fastclk_c_enable_35)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32189_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i32193_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n13805), 
         .Z(fastclk_c_enable_33)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32193_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i32187_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n13802), 
         .Z(fastclk_c_enable_36)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32187_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i32191_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n13803), 
         .Z(fastclk_c_enable_34)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32191_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i32195_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n13788), 
         .Z(fastclk_c_enable_32)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32195_3_lut_4_lut.init = 16'hd0f0;
    CCU2C _add_1_1284_add_4_11 (.A0(cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30470), .COUT(n30471), .S0(n54), .S1(n51));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_11.INJECT1_1 = "NO";
    LUT4 i32197_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n13806), 
         .Z(fastclk_c_enable_16)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32197_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_438 (.A(n1961), .B(n34354), .C(n13788), 
         .D(sda_in), .Z(n33438)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_438.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_439 (.A(n1961), .B(n34354), .C(n13802), 
         .D(sda_in), .Z(n33441)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_439.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_440 (.A(n1961), .B(n34354), .C(n27974), 
         .D(sda_in), .Z(n33440)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_440.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_441 (.A(n1961), .B(n34354), .C(n13806), 
         .D(sda_in), .Z(n33443)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_441.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_442 (.A(n1961), .B(n34354), .C(n13808), 
         .D(sda_in), .Z(n33439)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_442.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_443 (.A(n1961), .B(n34354), .C(n38349), 
         .D(sda_in), .Z(n33444)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_443.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_444 (.A(n1961), .B(n34354), .C(n13805), 
         .D(sda_in), .Z(n33442)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_444.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_445 (.A(n1961), .B(n34354), .C(n13803), 
         .D(sda_in), .Z(n33437)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_445.init = 16'h0200;
    LUT4 i32159_3_lut_4_lut (.A(n1961), .B(n34354), .C(n3572), .D(n38349), 
         .Z(fastclk_c_enable_5)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i32159_3_lut_4_lut.init = 16'hd0f0;
    LUT4 i1_3_lut_4_lut (.A(n1964), .B(n38324), .C(n1960), .D(n38338), 
         .Z(fastclk_c_enable_15)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_3_lut_4_lut.init = 16'hf2ff;
    LUT4 i1_3_lut_4_lut_adj_446 (.A(n1964), .B(n38324), .C(n453), .D(n2740), 
         .Z(n2741)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_3_lut_4_lut_adj_446.init = 16'hf200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_447 (.A(n1964), .B(n38324), .C(n3368), 
         .D(n1963), .Z(n10592)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_447.init = 16'h2f22;
    LUT4 i1_2_lut_4_lut (.A(n38347), .B(n38327), .C(n1965), .D(n33453), 
         .Z(n33454)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_4_lut.init = 16'h2000;
    LUT4 i1_3_lut_4_lut_adj_448 (.A(n36546), .B(n38328), .C(n33468), .D(rx_ready_N_322), 
         .Z(fastclk_c_enable_2)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_adj_448.init = 16'heefe;
    LUT4 mux_76_i2_3_lut_4_lut (.A(n38329), .B(n38347), .C(n2895), .D(bitidx[1]), 
         .Z(n487)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(181[34] 194[28])
    defparam mux_76_i2_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_76_i1_3_lut_4_lut (.A(n38329), .B(n38347), .C(n2895), .D(bitidx[0]), 
         .Z(n488)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(181[34] 194[28])
    defparam mux_76_i1_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_76_i3_3_lut_4_lut (.A(n38329), .B(n38347), .C(n2895), .D(bitidx[2]), 
         .Z(n486)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(181[34] 194[28])
    defparam mux_76_i3_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n38338), .B(n1968), .C(n38123), 
         .D(n1969), .Z(scl_t_N_310)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfffd;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n38338), .B(n36676), .C(n38330), .D(n1960), 
         .Z(fastclk_c_enable_45)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h5d55;
    LUT4 i1_3_lut_4_lut_4_lut_adj_449 (.A(n38338), .B(n36676), .C(n38330), 
         .D(n1960), .Z(fastclk_c_enable_91)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut_adj_449.init = 16'h5755;
    LUT4 i1149_4_lut_4_lut (.A(n38338), .B(n1961), .C(n34354), .D(n33454), 
         .Z(n3572)) /* synthesis lut_function=(!(A (B (C)+!B !(D)))) */ ;
    defparam i1149_4_lut_4_lut.init = 16'h7f5d;
    LUT4 i1_2_lut_rep_313_3_lut (.A(rx_ready_N_322), .B(n38336), .C(n1964), 
         .Z(n38318)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_313_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_450 (.A(rx_ready_N_322), .B(n38336), .C(n1964), 
         .Z(n81_adj_2261)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_3_lut_adj_450.init = 16'hefef;
    LUT4 i1_3_lut_4_lut_adj_451 (.A(n1960), .B(n38338), .C(rx_byte_idx[0]), 
         .D(rx_byte_idx[1]), .Z(n33457)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_3_lut_4_lut_adj_451.init = 16'h0880;
    CCU2C _add_1_1292_add_4_21 (.A0(gap[19]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[20]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30483), .COUT(n30484), .S0(n104), .S1(n101));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_452 (.A(cnt[6]), .B(n38337), .C(n38403), .D(rx_remaining[0]), 
         .Z(n30)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_4_lut_adj_452.init = 16'hfff7;
    LUT4 n31_bdd_2_lut_4_lut (.A(cnt[6]), .B(n38337), .C(n38403), .D(n38336), 
         .Z(n38121)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;
    defparam n31_bdd_2_lut_4_lut.init = 16'h00f7;
    LUT4 i709_2_lut_rep_306_4_lut (.A(cnt[6]), .B(n38337), .C(n38403), 
         .D(n38340), .Z(n38311)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i709_2_lut_rep_306_4_lut.init = 16'hf7ff;
    LUT4 i1_2_lut_4_lut_adj_453 (.A(cnt[6]), .B(n38337), .C(n38403), .D(n26), 
         .Z(n27)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_453.init = 16'h0800;
    LUT4 i1_2_lut_rep_307_4_lut (.A(cnt[6]), .B(n38337), .C(n38403), .D(rx_remaining[1]), 
         .Z(n38312)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_307_4_lut.init = 16'h0800;
    LUT4 i6643_2_lut_4_lut (.A(cnt[6]), .B(n38337), .C(n38403), .D(n1967), 
         .Z(n10583)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i6643_2_lut_4_lut.init = 16'hf700;
    CCU2C _add_1_1284_add_4_9 (.A0(cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30469), .COUT(n30470), .S0(n60_adj_2226), .S1(n57));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_9.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_9.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_9.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_25 (.A0(gap[23]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[24]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30485), .COUT(n30486), .S0(n92), .S1(n89));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_25.INJECT1_1 = "NO";
    CCU2C _add_1_1284_add_4_7 (.A0(cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30468), .COUT(n30469), .S0(n66_adj_2230), .S1(n63_adj_2223));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_7.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_7.INJECT1_1 = "NO";
    CCU2C _add_1_1284_add_4_5 (.A0(cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30467), .COUT(n30468), .S0(n72_adj_2227), .S1(n69_adj_2228));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_5.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_5.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_5.INJECT1_1 = "NO";
    CCU2C _add_1_1292_add_4_23 (.A0(gap[21]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[22]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30484), .COUT(n30485), .S0(n98), .S1(n95));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_23.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_23.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_23.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_321_4_lut (.A(n38350), .B(n38346), .C(cnt[6]), .D(n1964), 
         .Z(n38326)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_rep_321_4_lut.init = 16'h0400;
    LUT4 i22692_2_lut_rep_319_4_lut (.A(n38350), .B(n38346), .C(cnt[6]), 
         .D(rx_ready_N_322), .Z(n38324)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i22692_2_lut_rep_319_4_lut.init = 16'hfffb;
    LUT4 i1_3_lut_rep_322_4_lut (.A(n38346), .B(cnt[5]), .C(n38403), .D(cnt[6]), 
         .Z(n38327)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_3_lut_rep_322_4_lut.init = 16'hf7ff;
    LUT4 equal_314_i32_1_lut_rep_309_3_lut_4_lut (.A(n38346), .B(cnt[5]), 
         .C(n38403), .D(cnt[6]), .Z(fastclk_c_enable_47)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam equal_314_i32_1_lut_rep_309_3_lut_4_lut.init = 16'h0800;
    CCU2C _add_1_1284_add_4_3 (.A0(cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(cnt[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30466), .COUT(n30467), .S0(n78_adj_2220), .S1(n75_adj_2219));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_3.INIT0 = 16'haaa0;
    defparam _add_1_1284_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1284_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_3.INJECT1_1 = "NO";
    LUT4 i24462_2_lut_rep_333 (.A(rstn_c), .B(rst_N_5), .Z(n38338)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i24462_2_lut_rep_333.init = 16'h2222;
    LUT4 i1_2_lut_2_lut_3_lut (.A(rstn_c), .B(rst_N_5), .C(fastclk_c_enable_82), 
         .Z(fastclk_c_enable_83)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_2_lut_2_lut_3_lut.init = 16'hfdfd;
    CCU2C _add_1_1295_add_4_add_4_29 (.A0(n136), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30511), .S0(n3556));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_29.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_29.INIT1 = 16'h0000;
    defparam _add_1_1295_add_4_add_4_29.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_29.INJECT1_1 = "NO";
    LUT4 i24463_1_lut_rep_318_2_lut (.A(rstn_c), .B(rst_N_5), .Z(n38323)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i24463_1_lut_rep_318_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_305_3_lut_3_lut_4_lut (.A(rstn_c), .B(rst_N_5), .C(n1969), 
         .D(n1968), .Z(n38310)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_2_lut_rep_305_3_lut_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_323_3_lut (.A(rstn_c), .B(rst_N_5), .C(n2355), .Z(n38328)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_2_lut_rep_323_3_lut.init = 16'hfdfd;
    LUT4 i1_3_lut_3_lut_4_lut (.A(rstn_c), .B(rst_N_5), .C(n36620), .D(n34576), 
         .Z(fastclk_c_enable_31)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;
    defparam i1_3_lut_3_lut_4_lut.init = 16'hfddd;
    LUT4 i1_2_lut_rep_308_2_lut_3_lut (.A(rstn_c), .B(rst_N_5), .C(n1969), 
         .Z(n38313)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_2_lut_rep_308_2_lut_3_lut.init = 16'hfdfd;
    LUT4 i32171_3_lut_4_lut (.A(rstn_c), .B(rst_N_5), .C(n1969), .D(n38120), 
         .Z(sda_t_N_296)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i32171_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_2_lut_rep_320_3_lut (.A(rstn_c), .B(rst_N_5), .C(n1960), .Z(n38325)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_320_3_lut.init = 16'h2020;
    LUT4 i32166_2_lut_3_lut_4_lut (.A(rstn_c), .B(rst_N_5), .C(n38336), 
         .D(n1964), .Z(n33464)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i32166_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_2_lut_rep_315_3_lut_4_lut (.A(rstn_c), .B(rst_N_5), .C(n36546), 
         .D(n2355), .Z(fastclk_c_enable_3)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_2_lut_rep_315_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_4_lut_adj_454 (.A(n2960), .B(rx_ready), .C(n38348), 
         .D(reg_target[7]), .Z(reg_target_7__N_247[7])) /* synthesis lut_function=(A (D)+!A !(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_2_lut_4_lut_adj_454.init = 16'hba00;
    LUT4 i23883_2_lut_4_lut (.A(n2960), .B(rx_ready), .C(n38348), .D(reg_target[6]), 
         .Z(reg_target_7__N_247[6])) /* synthesis lut_function=(A (D)+!A !(B+!(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i23883_2_lut_4_lut.init = 16'hba00;
    IB rstn_pad (.I(rstn), .O(rstn_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(7[16:20])
    IB fastclk_pad (.I(fastclk), .O(fastclk_c));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(6[16:23])
    CCU2C _add_1_1295_add_4_add_4_27 (.A0(n58), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n136), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30510), .COUT(n30511), .S0(n66_adj_2216), .S1(n63_adj_2218));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_27.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_27.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_455 (.A(n38402), .B(n38350), .C(n38358), .D(n33370), 
         .Z(n20)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (D))) */ ;
    defparam i1_3_lut_4_lut_adj_455.init = 16'h20ff;
    LUT4 i1_2_lut_rep_337 (.A(n2353), .B(n38351), .Z(n38342)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_2_lut_rep_337.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_456 (.A(n2353), .B(n38351), .C(n2352), .Z(n13)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_2_lut_3_lut_adj_456.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_338 (.A(cnt[6]), .B(n15), .Z(n38343)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_338.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_457 (.A(cnt[6]), .B(n15), .C(n1876), 
         .D(n33370), .Z(n33465)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_457.init = 16'h0010;
    LUT4 i1_2_lut_rep_325_3_lut (.A(cnt[6]), .B(n15), .C(n33370), .Z(n38330)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_325_3_lut.init = 16'hfefe;
    LUT4 i31842_2_lut (.A(rx_byte_idx[0]), .B(rx_byte_idx[1]), .Z(n36676)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i31842_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_458 (.A(n36492), .B(n38403), .C(cnt[4]), .D(cnt[3]), 
         .Z(n33370)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_adj_458.init = 16'hfffe;
    LUT4 i1_2_lut_rep_299_3_lut_4_lut (.A(cnt[6]), .B(n15), .C(n1876), 
         .D(n33370), .Z(n38304)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_2_lut_rep_299_3_lut_4_lut.init = 16'hffef;
    CCU2C por_1137_add_4_17 (.A0(por[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30570), .S0(n70_adj_2215));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_17.INIT0 = 16'haaa0;
    defparam por_1137_add_4_17.INIT1 = 16'h0000;
    defparam por_1137_add_4_17.INJECT1_0 = "NO";
    defparam por_1137_add_4_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_459 (.A(cnt[5]), .B(cnt[2]), .Z(n36492)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_adj_459.init = 16'heeee;
    CCU2C por_1137_add_4_15 (.A0(por[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(por[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30569), .COUT(n30570), .S0(n72_adj_2213), .S1(n71_adj_2214));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_15.INIT0 = 16'haaa0;
    defparam por_1137_add_4_15.INIT1 = 16'haaa0;
    defparam por_1137_add_4_15.INJECT1_0 = "NO";
    defparam por_1137_add_4_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_339 (.A(tx_byte[0]), .B(n33384), .Z(n38344)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i1_2_lut_rep_339.init = 16'hdddd;
    LUT4 i994_3_lut_rep_324_4_lut (.A(tx_byte[0]), .B(n33384), .C(rx_ready_N_322), 
         .D(send_data_after_reg), .Z(n38329)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i994_3_lut_rep_324_4_lut.init = 16'h2f20;
    LUT4 i1_2_lut_3_lut_adj_460 (.A(tx_byte[0]), .B(n33384), .C(rx_ready_N_322), 
         .Z(n33453)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i1_2_lut_3_lut_adj_460.init = 16'h2020;
    LUT4 i1_2_lut_adj_461 (.A(n81_adj_2221), .B(n34), .Z(cnt_15__N_167[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_461.init = 16'h8888;
    CCU2C por_1137_add_4_13 (.A0(por[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(por[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30568), .COUT(n30569), .S0(n74_adj_2211), .S1(n73_adj_2212));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_13.INIT0 = 16'haaa0;
    defparam por_1137_add_4_13.INIT1 = 16'haaa0;
    defparam por_1137_add_4_13.INJECT1_0 = "NO";
    defparam por_1137_add_4_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_462 (.A(n15), .B(n34268), .C(n45_adj_2255), .D(n34606), 
         .Z(n34)) /* synthesis lut_function=(A (B+(D))+!A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_462.init = 16'hffdc;
    FD1P3AX por_1137__i15 (.D(n70_adj_2215), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i15.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_463 (.A(n15), .B(n38304), .C(n1969), .D(n103), 
         .Z(n34268)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(122[30] 129[28])
    defparam i1_4_lut_adj_463.init = 16'h0040;
    LUT4 i1_4_lut_adj_464 (.A(n1964), .B(n58_adj_2254), .C(n38402), .D(n55), 
         .Z(n45_adj_2255)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_464.init = 16'hceee;
    LUT4 i1_4_lut_adj_465 (.A(n15), .B(n38327), .C(n36696), .D(n103), 
         .Z(n34606)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_465.init = 16'h0004;
    LUT4 i1_4_lut_4_lut_adj_466 (.A(n38351), .B(rx_ready), .C(reg_target[0]), 
         .D(n2353), .Z(n3)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (D)+!B (C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_466.init = 16'h7400;
    LUT4 i1_3_lut_rep_331_4_lut (.A(n38402), .B(n15), .C(cnt[6]), .D(n38350), 
         .Z(n38336)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_3_lut_rep_331_4_lut.init = 16'hfffd;
    LUT4 i121_2_lut_rep_332_3_lut (.A(n38402), .B(n15), .C(cnt[5]), .Z(n38337)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i121_2_lut_rep_332_3_lut.init = 16'h2020;
    LUT4 i1_2_lut_rep_342 (.A(tx_byte[0]), .B(n33384), .Z(n38347)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i1_2_lut_rep_342.init = 16'heeee;
    LUT4 i22381_4_lut (.A(desired_read_len[1]), .B(n30), .C(n1960), .D(rx_remaining[1]), 
         .Z(rx_remaining_1__N_292[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i22381_4_lut.init = 16'hca0a;
    LUT4 i23445_2_lut_3_lut (.A(tx_byte[0]), .B(n33384), .C(reg_target[1]), 
         .Z(n452)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i23445_2_lut_3_lut.init = 16'h1010;
    LUT4 i31860_4_lut (.A(n1969), .B(n1963), .C(n1964), .D(n1959), .Z(n36696)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i31860_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_adj_467 (.A(cnt[6]), .B(n38402), .C(cnt[5]), .Z(n103)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_467.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_468 (.A(tx_byte[0]), .B(n33384), .C(reg_target[4]), 
         .Z(n449)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i1_2_lut_3_lut_adj_468.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(tx_byte[0]), .B(n33384), .C(n1965), 
         .D(n38327), .Z(n33468)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_4_lut_adj_469 (.A(n28124), .B(n34583), .C(n38324), .D(n1964), 
         .Z(fastclk_c_enable_82)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A ((C (D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_469.init = 16'h0c44;
    LUT4 i1_4_lut_adj_470 (.A(n38318), .B(n2740), .C(n38347), .D(n2651), 
         .Z(n34583)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_470.init = 16'hffbf;
    LUT4 i808_3_lut_4_lut (.A(tx_byte[0]), .B(n33384), .C(n38327), .D(n38329), 
         .Z(n2895)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i808_3_lut_4_lut.init = 16'hf0fe;
    LUT4 mux_69_i1_4_lut (.A(reg_target[0]), .B(n2651), .C(n38347), .D(write_data[0]), 
         .Z(n453)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(181[34] 194[28])
    defparam mux_69_i1_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_3_lut_adj_471 (.A(tx_byte[0]), .B(n33384), .C(reg_target[6]), 
         .Z(n447)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(178[29:55])
    defparam i1_2_lut_3_lut_adj_471.init = 16'h1010;
    LUT4 i688_2_lut (.A(send_data_after_reg), .B(rx_ready_N_322), .Z(n2651)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(189[34] 194[28])
    defparam i688_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_rep_334_4_lut (.A(n38406), .B(n2353), .C(rx_ready), 
         .D(n2960), .Z(n38339)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_3_lut_rep_334_4_lut.init = 16'hff0e;
    LUT4 i32174_4_lut (.A(n38338), .B(n38427), .C(n38324), .D(n1964), 
         .Z(n29256)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D))))) */ ;
    defparam i32174_4_lut.init = 16'h5f77;
    LUT4 i1_2_lut_3_lut_4_lut_adj_472 (.A(bitidx[0]), .B(n38401), .C(n1966), 
         .D(bitidx[3]), .Z(n36498)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(252[29:40])
    defparam i1_2_lut_3_lut_4_lut_adj_472.init = 16'hf0e0;
    LUT4 i1_2_lut_adj_473 (.A(n1969), .B(n1959), .Z(n3068)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_473.init = 16'heeee;
    LUT4 i1_4_lut_adj_474 (.A(rx_ready), .B(n38351), .C(n2354), .D(n2353), 
         .Z(n10610)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(38[9:17])
    defparam i1_4_lut_adj_474.init = 16'hf7a0;
    LUT4 i1_3_lut_adj_475 (.A(rx_ready), .B(n2355), .C(n2354), .Z(n10608)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(38[9:17])
    defparam i1_3_lut_adj_475.init = 16'hdcdc;
    LUT4 i6660_4_lut (.A(n1959), .B(rx_ready_N_322), .C(n38304), .D(n38326), 
         .Z(n10600)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i6660_4_lut.init = 16'heca0;
    LUT4 i6658_4_lut (.A(n1960), .B(n1961), .C(n38327), .D(n33398), 
         .Z(n10598)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i6658_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_476 (.A(bitidx[0]), .B(n13780), .C(n36672), .D(bitidx[1]), 
         .Z(n33398)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_476.init = 16'h0004;
    LUT4 i22940_2_lut_rep_303_3_lut_4_lut_4_lut (.A(bitidx[0]), .B(n38401), 
         .C(n38327), .D(bitidx[3]), .Z(n38308)) /* synthesis lut_function=(A+(B (C)+!B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(252[29:40])
    defparam i22940_2_lut_rep_303_3_lut_4_lut_4_lut.init = 16'hfafb;
    CCU2C _add_1_1295_add_4_add_4_25 (.A0(n60), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n59), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30509), .COUT(n30510), .S0(n72_adj_2217), .S1(n69_adj_2222));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_25.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_25.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_25.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_25.INJECT1_1 = "NO";
    LUT4 i31839_2_lut (.A(bitidx[2]), .B(bitidx[3]), .Z(n36672)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i31839_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_477 (.A(n38313), .B(n38343), .C(n66_adj_2231), .D(n56), 
         .Z(fastclk_c_enable_9)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(108[18] 361[12])
    defparam i1_4_lut_adj_477.init = 16'hfbfa;
    CCU2C por_1137_add_4_11 (.A0(por[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(por[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30567), .COUT(n30568), .S0(n76_adj_2209), .S1(n75_adj_2210));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_11.INIT0 = 16'haaa0;
    defparam por_1137_add_4_11.INIT1 = 16'haaa0;
    defparam por_1137_add_4_11.INJECT1_0 = "NO";
    defparam por_1137_add_4_11.INJECT1_1 = "NO";
    CCU2C por_1137_add_4_9 (.A0(por[7]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(por[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30566), 
          .COUT(n30567), .S0(n78_adj_2207), .S1(n77_adj_2208));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_9.INIT0 = 16'haaa0;
    defparam por_1137_add_4_9.INIT1 = 16'haaa0;
    defparam por_1137_add_4_9.INJECT1_0 = "NO";
    defparam por_1137_add_4_9.INJECT1_1 = "NO";
    LUT4 i70_3_lut (.A(n34062), .B(n3368), .C(n1963), .Z(n66_adj_2231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i70_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_478 (.A(n39283), .B(n34415), .C(n38341), .D(n33370), 
         .Z(n56)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i1_4_lut_adj_478.init = 16'h0ace;
    CCU2C por_1137_add_4_7 (.A0(por[5]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(por[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30565), 
          .COUT(n30566), .S0(n80_adj_2205), .S1(n79_adj_2206));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_7.INIT0 = 16'haaa0;
    defparam por_1137_add_4_7.INIT1 = 16'haaa0;
    defparam por_1137_add_4_7.INJECT1_0 = "NO";
    defparam por_1137_add_4_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_rep_346 (.A(rx_byte[7]), .B(n36576), .C(n36574), .D(rx_byte[2]), 
         .Z(n38351)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_rep_346.init = 16'hfffe;
    LUT4 i1_4_lut_adj_479 (.A(n38309), .B(n33453), .C(n7_adj_2260), .D(n33468), 
         .Z(n34410)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_479.init = 16'hfefa;
    LUT4 i13_4_lut (.A(n1961), .B(n1962), .C(n38327), .D(n38340), .Z(n7_adj_2260)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i13_4_lut.init = 16'hcac0;
    LUT4 i25_1_lut_rep_340_4_lut (.A(rx_byte[7]), .B(n36576), .C(n36574), 
         .D(rx_byte[2]), .Z(n38345)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i25_1_lut_rep_340_4_lut.init = 16'h0001;
    CCU2C por_1137_add_4_5 (.A0(por[3]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(por[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30564), 
          .COUT(n30565), .S0(n82_adj_2203), .S1(n81_adj_2204));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_5.INIT0 = 16'haaa0;
    defparam por_1137_add_4_5.INIT1 = 16'haaa0;
    defparam por_1137_add_4_5.INJECT1_0 = "NO";
    defparam por_1137_add_4_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_480 (.A(n34627), .B(n33469), .C(n1964), .D(n38336), 
         .Z(n34042)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_480.init = 16'hfeee;
    LUT4 i1_4_lut_adj_481 (.A(send_data_after_reg), .B(n33468), .C(n38344), 
         .D(rx_ready_N_322), .Z(n33469)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_481.init = 16'hc044;
    LUT4 i6648_4_lut (.A(n1965), .B(n1966), .C(n38327), .D(n33398), 
         .Z(n10588)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i6648_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_482 (.A(n10583), .B(n1968), .C(n38299), .D(n13780), 
         .Z(n36418)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_482.init = 16'hfefa;
    CCU2C por_1137_add_4_3 (.A0(por[1]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(por[2]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30563), 
          .COUT(n30564), .S0(n84), .S1(n83_adj_2202));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_3.INIT0 = 16'haaa0;
    defparam por_1137_add_4_3.INIT1 = 16'haaa0;
    defparam por_1137_add_4_3.INJECT1_0 = "NO";
    defparam por_1137_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_483 (.A(n38360), .B(n38359), .C(n36550), .D(n1959), 
         .Z(n34415)) /* synthesis lut_function=(A+(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_483.init = 16'hfafb;
    LUT4 i1_3_lut_adj_484 (.A(n1967), .B(n1963), .C(n1968), .Z(n36550)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_484.init = 16'hfefe;
    LUT4 i6642_4_lut (.A(n1968), .B(n1969), .C(n38327), .D(n33465), 
         .Z(n10582)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i6642_4_lut.init = 16'heca0;
    CCU2C por_1137_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(por[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30563), .S1(n85));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137_add_4_1.INIT0 = 16'h0000;
    defparam por_1137_add_4_1.INIT1 = 16'h555f;
    defparam por_1137_add_4_1.INJECT1_0 = "NO";
    defparam por_1137_add_4_1.INJECT1_1 = "NO";
    CCU2C _add_1_1295_add_4_add_4_23 (.A0(n62), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n61), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30508), .COUT(n30509), .S0(n78_adj_2224), .S1(n75_adj_2225));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_23.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_23.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_23.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_23.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_485 (.A(n1959), .B(n38310), .C(n36448), .D(n27), 
         .Z(fastclk_c_enable_10)) /* synthesis lut_function=(A (B)+!A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_485.init = 16'hdddc;
    LUT4 i1_4_lut_adj_486 (.A(n38343), .B(n26), .C(n20), .D(n23), .Z(n36448)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (C+(D))))) */ ;
    defparam i1_4_lut_adj_486.init = 16'h7350;
    CCU2C add_26226_32 (.A0(gap[31]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n30562), 
          .S1(n3368));
    defparam add_26226_32.INIT0 = 16'h555f;
    defparam add_26226_32.INIT1 = 16'h0000;
    defparam add_26226_32.INJECT1_0 = "NO";
    defparam add_26226_32.INJECT1_1 = "NO";
    PFUMX i32353 (.BLUT(n37740), .ALUT(n37739), .C0(bitidx[2]), .Z(n37741));
    CCU2C add_26226_30 (.A0(gap[29]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[30]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30561), 
          .COUT(n30562));
    defparam add_26226_30.INIT0 = 16'h555f;
    defparam add_26226_30.INIT1 = 16'h555f;
    defparam add_26226_30.INJECT1_0 = "NO";
    defparam add_26226_30.INJECT1_1 = "NO";
    CCU2C _add_1_1295_add_4_add_4_21 (.A0(n64), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n63), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30507), .COUT(n30508), .S0(n84_adj_2229), .S1(n81_adj_2232));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_21.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_21.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_21.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_21.INJECT1_1 = "NO";
    CCU2C _add_1_1295_add_4_add_4_19 (.A0(n66), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n65), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30506), .COUT(n30507), .S0(n90), .S1(n87));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_19.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_19.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_19.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_19.INJECT1_1 = "NO";
    CCU2C _add_1_1284_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cnt[0]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30466), .S1(n81_adj_2221));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(110[38:49])
    defparam _add_1_1284_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1284_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1284_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1284_add_4_1.INJECT1_1 = "NO";
    FD1P3IX rx_remaining__i1 (.D(rx_remaining_1__N_292[1]), .SP(fastclk_c_enable_15), 
            .CD(n38323), .CK(fastclk_c), .Q(rx_remaining[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_remaining__i1.GSR = "DISABLED";
    CCU2C add_26226_28 (.A0(gap[27]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[28]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30560), 
          .COUT(n30561));
    defparam add_26226_28.INIT0 = 16'h555f;
    defparam add_26226_28.INIT1 = 16'h555f;
    defparam add_26226_28.INJECT1_0 = "NO";
    defparam add_26226_28.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_487 (.A(n2960), .B(n3), .C(n13833), .D(reg_target[0]), 
         .Z(reg_target_7__N_247[0])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_4_lut_adj_487.init = 16'hfefc;
    CCU2C _add_1_1295_add_4_add_4_17 (.A0(n68), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n67), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30505), .COUT(n30506), .S0(n96), .S1(n93));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_17.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_17.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_17.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_488 (.A(n1967), .B(n1968), .C(n1962), .D(n1964), 
         .Z(n3070)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_488.init = 16'hfffe;
    LUT4 i1_2_lut_adj_489 (.A(n2349), .B(n2350), .Z(n2960)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_2_lut_adj_489.init = 16'heeee;
    LUT4 i32157_4_lut (.A(n29267), .B(n38338), .C(n3368), .D(n1963), 
         .Z(fastclk_c_enable_79)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C (D))))) */ ;
    defparam i32157_4_lut.init = 16'h3f77;
    LUT4 i25318_4_lut (.A(n3068), .B(n38324), .C(n1964), .D(n38330), 
         .Z(n29267)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i25318_4_lut.init = 16'hcfc5;
    LUT4 n31_bdd_3_lut_4_lut (.A(n1962), .B(n1967), .C(n38359), .D(n38327), 
         .Z(n38122)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam n31_bdd_3_lut_4_lut.init = 16'hf101;
    LUT4 i1_2_lut_3_lut_4_lut_adj_490 (.A(n1962), .B(n1967), .C(n1963), 
         .D(n3368), .Z(n23)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_490.init = 16'hfeee;
    LUT4 i1_2_lut_rep_353 (.A(n1960), .B(n1965), .Z(n38358)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_rep_353.init = 16'heeee;
    OB led_pad_0 (.I(led_c_0), .O(led[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(10[20:23])
    OB led_pad_1 (.I(led_c_1), .O(led[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(10[20:23])
    OB led_pad_2 (.I(led_c_2), .O(led[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(10[20:23])
    OB led_pad_3 (.I(led_c_3), .O(led[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(10[20:23])
    LUT4 i1_2_lut_rep_354 (.A(n1961), .B(n1966), .Z(n38359)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_rep_354.init = 16'heeee;
    LUT4 i22677_2_lut (.A(n161), .B(n32862), .Z(n2797)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i22677_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_491 (.A(n1961), .B(n1966), .C(n1965), 
         .D(n1960), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_3_lut_4_lut_adj_491.init = 16'hfffe;
    LUT4 i1_2_lut_rep_355 (.A(n1969), .B(n1964), .Z(n38360)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_rep_355.init = 16'heeee;
    LUT4 i1_4_lut_4_lut_adj_492 (.A(n1969), .B(n1964), .C(n1967), .D(n1968), 
         .Z(n34062)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_4_lut_adj_492.init = 16'h0302;
    FD1P3IX rx_byte__i1 (.D(n33443), .SP(fastclk_c_enable_16), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_493 (.A(bitidx[0]), .B(bitidx[2]), .C(bitidx[1]), 
         .Z(n13808)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_adj_493.init = 16'hf7f7;
    LUT4 i24024_2_lut_3_lut (.A(bitidx[0]), .B(bitidx[2]), .C(bitidx[1]), 
         .Z(n27974)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i24024_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_494 (.A(bitidx[0]), .B(bitidx[2]), .C(bitidx[1]), 
         .Z(n13803)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_3_lut_adj_494.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_495 (.A(bitidx[0]), .B(bitidx[2]), .C(bitidx[1]), 
         .Z(n13802)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_3_lut_adj_495.init = 16'hbfbf;
    LUT4 i1_2_lut_3_lut_adj_496 (.A(bitidx[2]), .B(bitidx[1]), .C(bitidx[0]), 
         .Z(n13788)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_3_lut_adj_496.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_497 (.A(bitidx[2]), .B(bitidx[1]), .C(bitidx[0]), 
         .Z(n13805)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_3_lut_adj_497.init = 16'hbfbf;
    CCU2C _add_1_1295_add_4_add_4_15 (.A0(n70), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n69), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30504), .COUT(n30505), .S0(n102), .S1(n99));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_15.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_15.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_15.INJECT1_1 = "NO";
    CCU2C _add_1_1295_add_4_add_4_13 (.A0(n72), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n71), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30503), .COUT(n30504), .S0(n108), .S1(n105));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_13.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_13.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_13.INJECT1_1 = "NO";
    FD1P3AX por_1137__i14 (.D(n71_adj_2214), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i14.GSR = "DISABLED";
    FD1P3AX por_1137__i13 (.D(n72_adj_2213), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i13.GSR = "DISABLED";
    FD1P3AX por_1137__i12 (.D(n73_adj_2212), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i12.GSR = "DISABLED";
    FD1P3AX por_1137__i11 (.D(n74_adj_2211), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i11.GSR = "DISABLED";
    FD1P3AX por_1137__i10 (.D(n75_adj_2210), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i10.GSR = "DISABLED";
    FD1P3AX por_1137__i9 (.D(n76_adj_2209), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i9.GSR = "DISABLED";
    FD1P3AX por_1137__i8 (.D(n77_adj_2208), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i8.GSR = "DISABLED";
    FD1P3AX por_1137__i7 (.D(n78_adj_2207), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i7.GSR = "DISABLED";
    FD1P3AX por_1137__i6 (.D(n79_adj_2206), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i6.GSR = "DISABLED";
    FD1P3AX por_1137__i5 (.D(n80_adj_2205), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i5.GSR = "DISABLED";
    FD1P3AX por_1137__i4 (.D(n81_adj_2204), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i4.GSR = "DISABLED";
    FD1P3AX por_1137__i3 (.D(n82_adj_2203), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i3.GSR = "DISABLED";
    FD1P3AX por_1137__i2 (.D(n83_adj_2202), .SP(rst_N_5), .CK(fastclk_c), 
            .Q(por[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i2.GSR = "DISABLED";
    FD1P3AX por_1137__i1 (.D(n84), .SP(rst_N_5), .CK(fastclk_c), .Q(por[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(18[37:48])
    defparam por_1137__i1.GSR = "DISABLED";
    FD1P3IX distance__i15 (.D(msb[7]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i15.GSR = "DISABLED";
    FD1P3IX distance__i14 (.D(msb[6]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i14.GSR = "DISABLED";
    FD1P3IX distance__i13 (.D(msb[5]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i13.GSR = "DISABLED";
    FD1P3IX distance__i12 (.D(msb[4]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i12.GSR = "DISABLED";
    FD1P3IX distance__i11 (.D(msb[3]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i11.GSR = "DISABLED";
    FD1P3IX distance__i10 (.D(msb[2]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i10.GSR = "DISABLED";
    FD1P3IX distance__i9 (.D(msb[1]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i9.GSR = "DISABLED";
    FD1P3IX distance__i8 (.D(msb[0]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i8.GSR = "DISABLED";
    FD1P3IX distance__i7 (.D(lsb[7]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i7.GSR = "DISABLED";
    FD1P3IX distance__i6 (.D(lsb[6]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i6.GSR = "DISABLED";
    FD1P3IX distance__i5 (.D(lsb[5]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i5.GSR = "DISABLED";
    FD1P3IX distance__i4 (.D(lsb[4]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i4.GSR = "DISABLED";
    FD1P3IX distance__i3 (.D(lsb[3]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i3.GSR = "DISABLED";
    FD1P3IX distance__i2 (.D(lsb[2]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i2.GSR = "DISABLED";
    FD1P3IX distance__i1 (.D(lsb[1]), .SP(fastclk_c_enable_31), .CD(n38323), 
            .CK(fastclk_c), .Q(distance[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam distance__i1.GSR = "DISABLED";
    FD1S3IX seq_state_FSM_i6 (.D(n36620), .CK(fastclk_c), .CD(n38323), 
            .Q(n2349));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam seq_state_FSM_i6.GSR = "DISABLED";
    FD1P3IX rx_byte__i2 (.D(n33438), .SP(fastclk_c_enable_32), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i2.GSR = "DISABLED";
    FD1P3IX rx_byte__i3 (.D(n33442), .SP(fastclk_c_enable_33), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i3.GSR = "DISABLED";
    FD1P3IX rx_byte__i4 (.D(n33437), .SP(fastclk_c_enable_34), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i4.GSR = "DISABLED";
    FD1P3IX rx_byte__i5 (.D(n33439), .SP(fastclk_c_enable_35), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i5.GSR = "DISABLED";
    FD1P3IX rx_byte__i6 (.D(n33441), .SP(fastclk_c_enable_36), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i6.GSR = "DISABLED";
    FD1P3IX rx_byte__i7 (.D(n33440), .SP(fastclk_c_enable_37), .CD(n38323), 
            .CK(fastclk_c), .Q(rx_byte[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte__i7.GSR = "DISABLED";
    FD1P3JX tx_byte_i1 (.D(n452), .SP(fastclk_c_enable_83), .PD(n29256), 
            .CK(fastclk_c), .Q(tx_byte[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i1.GSR = "DISABLED";
    FD1S3IX seq_state_FSM_i5 (.D(n10614), .CK(fastclk_c), .CD(n38323), 
            .Q(n2350));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam seq_state_FSM_i5.GSR = "DISABLED";
    FD1P3IX seq_state_FSM_i4 (.D(n38342), .SP(rx_ready), .CD(n38323), 
            .CK(fastclk_c), .Q(n2352));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam seq_state_FSM_i4.GSR = "DISABLED";
    FD1S3IX seq_state_FSM_i3 (.D(n10610), .CK(fastclk_c), .CD(n38323), 
            .Q(n2353));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam seq_state_FSM_i3.GSR = "DISABLED";
    FD1S3IX seq_state_FSM_i2 (.D(n10608), .CK(fastclk_c), .CD(n38323), 
            .Q(n2354));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam seq_state_FSM_i2.GSR = "DISABLED";
    FD1P3IX lsb__i7 (.D(rx_byte[7]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i7.GSR = "DISABLED";
    FD1P3IX lsb__i6 (.D(rx_byte[6]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i6.GSR = "DISABLED";
    FD1P3IX lsb__i5 (.D(rx_byte[5]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i5.GSR = "DISABLED";
    FD1P3IX lsb__i4 (.D(rx_byte[4]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i4.GSR = "DISABLED";
    FD1P3IX lsb__i3 (.D(rx_byte[3]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i3.GSR = "DISABLED";
    FD1P3IX lsb__i2 (.D(rx_byte[2]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i2.GSR = "DISABLED";
    FD1P3IX lsb__i1 (.D(rx_byte[1]), .SP(fastclk_c_enable_45), .CD(n38323), 
            .CK(fastclk_c), .Q(lsb[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam lsb__i1.GSR = "DISABLED";
    FD1S3IX state_FSM_i11 (.D(n10600), .CK(fastclk_c), .CD(n38323), .Q(n1959));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i11.GSR = "DISABLED";
    FD1S3IX state_FSM_i10 (.D(n10598), .CK(fastclk_c), .CD(n38323), .Q(n1960));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i10.GSR = "DISABLED";
    FD1P3IX state_FSM_i9 (.D(n1962), .SP(fastclk_c_enable_47), .CD(n38323), 
            .CK(fastclk_c), .Q(n1961));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i9.GSR = "DISABLED";
    FD1S3IX state_FSM_i8 (.D(n34410), .CK(fastclk_c), .CD(n38323), .Q(n1962));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i8.GSR = "DISABLED";
    FD1S3IX state_FSM_i7 (.D(n10592), .CK(fastclk_c), .CD(n38323), .Q(n1963));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i7.GSR = "DISABLED";
    FD1S3IX state_FSM_i6 (.D(n34042), .CK(fastclk_c), .CD(n38323), .Q(n1964));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i6.GSR = "DISABLED";
    FD1S3IX state_FSM_i5 (.D(n10588), .CK(fastclk_c), .CD(n38323), .Q(n1965));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i5.GSR = "DISABLED";
    FD1P3IX state_FSM_i4 (.D(n1967), .SP(fastclk_c_enable_47), .CD(n38323), 
            .CK(fastclk_c), .Q(n1966));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i4.GSR = "DISABLED";
    FD1S3IX state_FSM_i3 (.D(n34303), .CK(fastclk_c), .CD(n38323), .Q(n1967));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n10582), .CK(fastclk_c), .CD(n38323), .Q(n1968));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1P3IX gap__i31 (.D(n2828), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i31.GSR = "DISABLED";
    CCU2C _add_1_1295_add_4_add_4_11 (.A0(n74), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n73), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30502), .COUT(n30503), .S0(n114), .S1(n111));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_11.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_11.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_11.INJECT1_1 = "NO";
    CCU2C add_26226_26 (.A0(gap[25]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[26]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30559), 
          .COUT(n30560));
    defparam add_26226_26.INIT0 = 16'h555f;
    defparam add_26226_26.INIT1 = 16'h555f;
    defparam add_26226_26.INJECT1_0 = "NO";
    defparam add_26226_26.INJECT1_1 = "NO";
    LUT4 i1_4_lut_then_4_lut (.A(n3070), .B(n1960), .C(n3068), .D(n1963), 
         .Z(n38420)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_then_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_else_4_lut (.A(n3368), .B(n3068), .C(n38304), .D(n1963), 
         .Z(n38419)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_else_4_lut.init = 16'hae0c;
    LUT4 i1_4_lut_then_3_lut (.A(n1876), .B(n1963), .C(n3368), .Z(n38423)) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_then_3_lut.init = 16'ha2a2;
    LUT4 i1_4_lut_else_3_lut (.A(n1876), .B(n1963), .C(n3368), .D(n1964), 
         .Z(n38422)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_else_3_lut.init = 16'hb3a2;
    LUT4 i28_4_lut_then_4_lut (.A(n38327), .B(n1964), .C(n38336), .D(rx_ready_N_322), 
         .Z(n38426)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i28_4_lut_then_4_lut.init = 16'hbbbf;
    LUT4 i28_4_lut_else_4_lut (.A(n38343), .B(n33370), .C(n3068), .D(n1876), 
         .Z(n38425)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i28_4_lut_else_4_lut.init = 16'hefff;
    LUT4 n5_bdd_3_lut_32486_then_3_lut (.A(tx_byte[6]), .B(tx_byte[7]), 
         .C(bitidx[0]), .Z(n38429)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam n5_bdd_3_lut_32486_then_3_lut.init = 16'h3535;
    LUT4 n5_bdd_3_lut_32486_else_3_lut (.A(tx_byte[3]), .B(tx_byte[2]), 
         .C(bitidx[0]), .Z(n38428)) /* synthesis lut_function=(!(A (B+(C))+!A !((C)+!B))) */ ;
    defparam n5_bdd_3_lut_32486_else_3_lut.init = 16'h5353;
    FD1P3IX gap__i30 (.D(n2827), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i30.GSR = "DISABLED";
    FD1P3IX gap__i29 (.D(n2826), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i29.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_498 (.A(n36456), .B(bitidx[0]), .C(n38359), .D(n38311), 
         .Z(bitidx_3__N_195[0])) /* synthesis lut_function=(A+(B (C (D))+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_498.init = 16'heaba;
    FD1P3IX gap__i28 (.D(n2825), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i28.GSR = "DISABLED";
    FD1P3IX gap__i27 (.D(n2824), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i27.GSR = "DISABLED";
    FD1P3IX gap__i26 (.D(n2823), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i26.GSR = "DISABLED";
    FD1P3IX gap__i25 (.D(n2822), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i25.GSR = "DISABLED";
    LUT4 n29978_bdd_4_lut (.A(n38328), .B(n2354), .C(rx_ready), .D(n2352), 
         .Z(n14113)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam n29978_bdd_4_lut.init = 16'hfaea;
    FD1P3IX gap__i24 (.D(n2821), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i24.GSR = "DISABLED";
    FD1P3IX gap__i23 (.D(n2820), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i23.GSR = "DISABLED";
    FD1P3IX gap__i22 (.D(n2819), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i22.GSR = "DISABLED";
    FD1P3IX gap__i21 (.D(n2818), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i21.GSR = "DISABLED";
    FD1P3IX gap__i20 (.D(n2817), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i20.GSR = "DISABLED";
    FD1P3IX gap__i19 (.D(n2816), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i19.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_499 (.A(n488), .B(n38309), .C(n38421), .D(n1965), 
         .Z(n36456)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_499.init = 16'hfefc;
    LUT4 n37741_bdd_3_lut (.A(n1960), .B(rx_remaining[1]), .C(n1968), 
         .Z(n38117)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam n37741_bdd_3_lut.init = 16'hf8f8;
    LUT4 n37741_bdd_3_lut_32480 (.A(n37741), .B(n38430), .C(bitidx[1]), 
         .Z(n38116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n37741_bdd_3_lut_32480.init = 16'hcaca;
    LUT4 i433_2_lut_rep_294 (.A(n3368), .B(n1963), .Z(n38299)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i433_2_lut_rep_294.init = 16'h8888;
    LUT4 n38118_bdd_3_lut (.A(n38118), .B(n38336), .C(n1964), .Z(n38119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38118_bdd_3_lut.init = 16'hcaca;
    LUT4 i24173_3_lut_4_lut (.A(n38304), .B(n3068), .C(n1965), .D(n38327), 
         .Z(n28124)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i24173_3_lut_4_lut.init = 16'hfb0b;
    FD1P3IX gap__i18 (.D(n2815), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i18.GSR = "DISABLED";
    FD1P3IX gap__i17 (.D(n2814), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i17.GSR = "DISABLED";
    FD1P3IX gap__i16 (.D(n2813), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i16.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_297 (.A(n1963), .B(n3368), .Z(n38302)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_rep_297.init = 16'h2222;
    FD1P3IX gap__i15 (.D(n2812), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i15.GSR = "DISABLED";
    LUT4 n38119_bdd_3_lut (.A(n38119), .B(n3368), .C(n1963), .Z(n38120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38119_bdd_3_lut.init = 16'hcaca;
    FD1P3IX gap__i14 (.D(n2811), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i14.GSR = "DISABLED";
    FD1P3IX gap__i13 (.D(n2810), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i13.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_500 (.A(n1963), .B(n3368), .C(n1959), .D(n103), 
         .Z(n58_adj_2254)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_3_lut_4_lut_adj_500.init = 16'h00f2;
    FD1P3JX tx_byte_i4 (.D(n449), .SP(fastclk_c_enable_83), .PD(n29256), 
            .CK(fastclk_c), .Q(tx_byte[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i4.GSR = "DISABLED";
    FD1P3IX gap__i12 (.D(n2809), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i12.GSR = "DISABLED";
    FD1P3IX gap__i11 (.D(n2808), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i11.GSR = "DISABLED";
    FD1P3IX gap__i10 (.D(n2807), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i10.GSR = "DISABLED";
    FD1P3IX gap__i9 (.D(n2806), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i9.GSR = "DISABLED";
    FD1P3IX gap__i8 (.D(n2805), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i8.GSR = "DISABLED";
    LUT4 select_853_Select_1_i6_3_lut_4_lut (.A(n38330), .B(n1876), .C(n3068), 
         .D(bitidx[1]), .Z(n6_adj_2259)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam select_853_Select_1_i6_3_lut_4_lut.init = 16'hf040;
    FD1P3IX gap__i7 (.D(n2804), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i7.GSR = "DISABLED";
    LUT4 select_853_Select_2_i6_3_lut_4_lut (.A(n38330), .B(n1876), .C(n3068), 
         .D(bitidx[2]), .Z(n6)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;
    defparam select_853_Select_2_i6_3_lut_4_lut.init = 16'hf040;
    LUT4 n1964_bdd_2_lut (.A(n1964), .B(n1963), .Z(n39283)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n1964_bdd_2_lut.init = 16'h2222;
    FD1P3IX gap__i6 (.D(n2803), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i6.GSR = "DISABLED";
    CCU2C _add_1_1295_add_4_add_4_9 (.A0(n76), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n75), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30501), .COUT(n30502), .S0(n120), .S1(n117));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_9.INJECT1_1 = "NO";
    FD1P3IX gap__i5 (.D(n2802), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i5.GSR = "DISABLED";
    FD1P3IX gap__i4 (.D(n2801), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i4.GSR = "DISABLED";
    FD1P3IX gap__i3 (.D(n2800), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i3.GSR = "DISABLED";
    FD1P3IX gap__i2 (.D(n2799), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i2.GSR = "DISABLED";
    FD1P3IX gap__i1 (.D(n2798), .SP(fastclk_c_enable_79), .CD(n38323), 
            .CK(fastclk_c), .Q(gap[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam gap__i1.GSR = "DISABLED";
    FD1S3JX reg_target_i7 (.D(reg_target_7__N_247[7]), .CK(fastclk_c), .PD(n38323), 
            .Q(reg_target[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i7.GSR = "DISABLED";
    FD1S3JX reg_target_i6 (.D(reg_target_7__N_247[6]), .CK(fastclk_c), .PD(n38323), 
            .Q(reg_target[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i6.GSR = "DISABLED";
    FD1S3IX reg_target_i4 (.D(reg_target_7__N_247[4]), .CK(fastclk_c), .CD(n38323), 
            .Q(reg_target[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i4.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_501 (.A(desired_read_len[1]), .B(desired_read_len[0]), 
         .Z(n28)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_adj_501.init = 16'hdddd;
    FD1S3IX reg_target_i3 (.D(reg_target_7__N_247[3]), .CK(fastclk_c), .CD(n38323), 
            .Q(reg_target[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i3.GSR = "DISABLED";
    FD1S3IX reg_target_i2 (.D(reg_target_7__N_247[2]), .CK(fastclk_c), .CD(n38323), 
            .Q(reg_target[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i2.GSR = "DISABLED";
    FD1S3JX reg_target_i1 (.D(reg_target_7__N_247[1]), .CK(fastclk_c), .PD(n38323), 
            .Q(reg_target[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam reg_target_i1.GSR = "DISABLED";
    FD1P3IX tx_byte_i7 (.D(n2748), .SP(fastclk_c_enable_82), .CD(n38323), 
            .CK(fastclk_c), .Q(tx_byte[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i7.GSR = "DISABLED";
    CCU2C _add_1_1292_add_4_27 (.A0(gap[25]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(gap[26]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30486), .COUT(n30487), .S0(n86), .S1(n83_adj_2238));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(288[52:63])
    defparam _add_1_1292_add_4_27.INIT0 = 16'haaa0;
    defparam _add_1_1292_add_4_27.INIT1 = 16'haaa0;
    defparam _add_1_1292_add_4_27.INJECT1_0 = "NO";
    defparam _add_1_1292_add_4_27.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_502 (.A(rx_byte[3]), .B(rx_byte[5]), .C(rx_byte[0]), 
         .D(rx_byte[4]), .Z(n36576)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_502.init = 16'hfffe;
    LUT4 i1_2_lut_adj_503 (.A(rx_byte[6]), .B(rx_byte[1]), .Z(n36574)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_503.init = 16'heeee;
    FD1P3IX tx_byte_i3 (.D(n2744), .SP(fastclk_c_enable_82), .CD(n38323), 
            .CK(fastclk_c), .Q(tx_byte[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i3.GSR = "DISABLED";
    FD1P3IX tx_byte_i2 (.D(n2743), .SP(fastclk_c_enable_82), .CD(n38323), 
            .CK(fastclk_c), .Q(tx_byte[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i2.GSR = "DISABLED";
    LUT4 i32181_4_lut (.A(n36528), .B(n36540), .C(n36538), .D(n36522), 
         .Z(rst_N_5)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i32181_4_lut.init = 16'h7fff;
    LUT4 i1_2_lut_adj_504 (.A(por[3]), .B(por[9]), .Z(n36528)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_504.init = 16'h8888;
    LUT4 i1_4_lut_adj_505 (.A(por[14]), .B(n36536), .C(n36530), .D(por[13]), 
         .Z(n36540)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_505.init = 16'h8000;
    CCU2C add_26226_24 (.A0(gap[23]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[24]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30558), 
          .COUT(n30559));
    defparam add_26226_24.INIT0 = 16'h555f;
    defparam add_26226_24.INIT1 = 16'h555f;
    defparam add_26226_24.INJECT1_0 = "NO";
    defparam add_26226_24.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_506 (.A(por[15]), .B(por[8]), .C(por[1]), .D(por[6]), 
         .Z(n36538)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_506.init = 16'h8000;
    LUT4 i1_2_lut_adj_507 (.A(por[2]), .B(por[4]), .Z(n36522)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_507.init = 16'h8888;
    FD1S3IX cnt__i15 (.D(cnt_15__N_167[15]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[15])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i15.GSR = "DISABLED";
    FD1S3IX cnt__i14 (.D(cnt_15__N_167[14]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[14])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i14.GSR = "DISABLED";
    FD1S3IX cnt__i13 (.D(cnt_15__N_167[13]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[13])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i13.GSR = "DISABLED";
    FD1S3IX cnt__i12 (.D(cnt_15__N_167[12]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[12])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i12.GSR = "DISABLED";
    FD1S3IX cnt__i11 (.D(cnt_15__N_167[11]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[11])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i11.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_508 (.A(por[10]), .B(por[7]), .C(por[0]), .D(por[11]), 
         .Z(n36536)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_508.init = 16'h8000;
    LUT4 i1_2_lut_adj_509 (.A(por[5]), .B(por[12]), .Z(n36530)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_509.init = 16'h8888;
    FD1S3IX cnt__i10 (.D(cnt_15__N_167[10]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[10])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i10.GSR = "DISABLED";
    FD1S3IX cnt__i9 (.D(cnt_15__N_167[9]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[9])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i9.GSR = "DISABLED";
    FD1S3IX cnt__i8 (.D(cnt_15__N_167[8]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[8])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i8.GSR = "DISABLED";
    FD1S3IX cnt__i7 (.D(cnt_15__N_167[7]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[7])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i7.GSR = "DISABLED";
    FD1S3IX cnt__i6 (.D(cnt_15__N_167[6]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[6])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i6.GSR = "DISABLED";
    FD1S3IX cnt__i5 (.D(cnt_15__N_167[5]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[5])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i5.GSR = "DISABLED";
    CCU2C add_26226_22 (.A0(gap[21]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[22]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30557), 
          .COUT(n30558));
    defparam add_26226_22.INIT0 = 16'h555f;
    defparam add_26226_22.INIT1 = 16'h555f;
    defparam add_26226_22.INJECT1_0 = "NO";
    defparam add_26226_22.INJECT1_1 = "NO";
    FD1S3IX cnt__i4 (.D(cnt_15__N_167[4]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[4])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i4.GSR = "DISABLED";
    FD1S3IX cnt__i3 (.D(cnt_15__N_167[3]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[3])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i3.GSR = "DISABLED";
    FD1S3IX cnt__i2 (.D(cnt_15__N_167[2]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[2])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i2.GSR = "DISABLED";
    FD1S3IX cnt__i1 (.D(cnt_15__N_167[1]), .CK(fastclk_c), .CD(n38323), 
            .Q(cnt[1])) /* synthesis lse_init_val=0 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam cnt__i1.GSR = "DISABLED";
    CCU2C _add_1_1295_add_4_add_4_7 (.A0(n78), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n77), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30500), .COUT(n30501), .S0(n126), .S1(n123));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_7.INIT0 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_7.INIT1 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_7.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_7.INJECT1_1 = "NO";
    FD1P3JX tx_byte_i6 (.D(n447), .SP(fastclk_c_enable_83), .PD(n29256), 
            .CK(fastclk_c), .Q(tx_byte[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam tx_byte_i6.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_510 (.A(n38338), .B(n38404), .C(n2355), .D(n38405), 
         .Z(n3638)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(16[16:44])
    defparam i1_4_lut_adj_510.init = 16'ha0a8;
    LUT4 i1_4_lut_adj_511 (.A(n2), .B(n36480), .C(n36474), .D(n3_adj_2257), 
         .Z(rx_ready_N_322)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam i1_4_lut_adj_511.init = 16'hfffe;
    LUT4 tx_byte_7__I_0_307_i2_2_lut (.A(tx_byte[1]), .B(reg_target[1]), 
         .Z(n2)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam tx_byte_7__I_0_307_i2_2_lut.init = 16'h6666;
    LUT4 i1_4_lut_adj_512 (.A(n5_adj_2256), .B(n1), .C(tx_byte[3]), .D(reg_target[3]), 
         .Z(n36480)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(205[29:50])
    defparam i1_4_lut_adj_512.init = 16'heffe;
    CCU2C add_26226_20 (.A0(gap[19]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[20]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30556), 
          .COUT(n30557));
    defparam add_26226_20.INIT0 = 16'h555f;
    defparam add_26226_20.INIT1 = 16'h555f;
    defparam add_26226_20.INJECT1_0 = "NO";
    defparam add_26226_20.INJECT1_1 = "NO";
    CCU2C _add_1_1295_add_4_add_4_5 (.A0(n80), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n79), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30499), .COUT(n30500), .S0(n132), .S1(n129));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_5.INIT0 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_5.INIT1 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_5.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_5.INJECT1_1 = "NO";
    CCU2C add_26226_18 (.A0(gap[17]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[18]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30555), 
          .COUT(n30556));
    defparam add_26226_18.INIT0 = 16'h555f;
    defparam add_26226_18.INIT1 = 16'h555f;
    defparam add_26226_18.INJECT1_0 = "NO";
    defparam add_26226_18.INJECT1_1 = "NO";
    FD1P3IX msb__i7 (.D(rx_byte[7]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i7.GSR = "DISABLED";
    LUT4 tx_byte_0__bdd_2_lut_32991 (.A(tx_byte[4]), .B(bitidx[0]), .Z(n37739)) /* synthesis lut_function=((B)+!A) */ ;
    defparam tx_byte_0__bdd_2_lut_32991.init = 16'hdddd;
    CCU2C _add_1_1295_add_4_add_4_3 (.A0(n82), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n81), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30498), .COUT(n30499), .S0(n138), .S1(n135));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_3.INIT0 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_3.INIT1 = 16'haaa0;
    defparam _add_1_1295_add_4_add_4_3.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_3.INJECT1_1 = "NO";
    CCU2C add_26226_16 (.A0(gap[15]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30554), 
          .COUT(n30555));
    defparam add_26226_16.INIT0 = 16'h555f;
    defparam add_26226_16.INIT1 = 16'h555f;
    defparam add_26226_16.INJECT1_0 = "NO";
    defparam add_26226_16.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_513 (.A(n36428), .B(bitidx[1]), .C(n38359), .D(n38308), 
         .Z(bitidx_3__N_195[1])) /* synthesis lut_function=(A+(B (C (D))+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_513.init = 16'heaba;
    LUT4 i1_4_lut_adj_514 (.A(bitidx[1]), .B(n36426), .C(n1960), .D(n38312), 
         .Z(n36428)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_514.init = 16'hfcec;
    CCU2C add_26226_14 (.A0(gap[13]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30553), 
          .COUT(n30554));
    defparam add_26226_14.INIT0 = 16'h555f;
    defparam add_26226_14.INIT1 = 16'h555f;
    defparam add_26226_14.INJECT1_0 = "NO";
    defparam add_26226_14.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_515 (.A(n487), .B(n6_adj_2259), .C(n1965), .D(n36422), 
         .Z(n36426)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_515.init = 16'hffec;
    LUT4 i1_4_lut_adj_516 (.A(bitidx[1]), .B(n3070), .C(n1963), .D(n3368), 
         .Z(n36422)) /* synthesis lut_function=(A (B+(C))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_516.init = 16'hf8a8;
    LUT4 i1_4_lut_adj_517 (.A(n36412), .B(bitidx[2]), .C(n38359), .D(n33483), 
         .Z(bitidx_3__N_195[2])) /* synthesis lut_function=(A+(B (C (D))+!B !((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_517.init = 16'heaba;
    CCU2C _add_1_1295_add_4_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n83), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30498), .S1(n141));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:38])
    defparam _add_1_1295_add_4_add_4_1.INIT0 = 16'h0000;
    defparam _add_1_1295_add_4_add_4_1.INIT1 = 16'h555f;
    defparam _add_1_1295_add_4_add_4_1.INJECT1_0 = "NO";
    defparam _add_1_1295_add_4_add_4_1.INJECT1_1 = "NO";
    CCU2C add_26226_12 (.A0(gap[11]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30552), 
          .COUT(n30553));
    defparam add_26226_12.INIT0 = 16'h555f;
    defparam add_26226_12.INIT1 = 16'h555f;
    defparam add_26226_12.INJECT1_0 = "NO";
    defparam add_26226_12.INJECT1_1 = "NO";
    FD1P3AX rx_byte_idx__i1 (.D(n33457), .SP(fastclk_c_enable_85), .CK(fastclk_c), 
            .Q(rx_byte_idx[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam rx_byte_idx__i1.GSR = "DISABLED";
    FD1P3IX msb__i6 (.D(rx_byte[6]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i6.GSR = "DISABLED";
    FD1P3IX msb__i5 (.D(rx_byte[5]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i5.GSR = "DISABLED";
    FD1P3IX msb__i4 (.D(rx_byte[4]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i4.GSR = "DISABLED";
    FD1P3IX msb__i3 (.D(rx_byte[3]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i3.GSR = "DISABLED";
    FD1P3IX msb__i2 (.D(rx_byte[2]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i2.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_518 (.A(n1960), .B(n36410), .C(bitidx[2]), .D(n38312), 
         .Z(n36412)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_518.init = 16'heeec;
    FD1P3IX msb__i1 (.D(rx_byte[1]), .SP(fastclk_c_enable_91), .CD(n38323), 
            .CK(fastclk_c), .Q(msb[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam msb__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_396 (.A(bitidx[1]), .B(bitidx[2]), .Z(n38401)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_rep_396.init = 16'heeee;
    LUT4 i1_2_lut_rep_344_3_lut (.A(bitidx[1]), .B(bitidx[2]), .C(bitidx[0]), 
         .Z(n38349)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_rep_344_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_519 (.A(bitidx[1]), .B(bitidx[2]), .C(bitidx[0]), 
         .Z(n13806)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_3_lut_adj_519.init = 16'hefef;
    LUT4 i1_2_lut_rep_335_3_lut_4_lut (.A(bitidx[1]), .B(bitidx[2]), .C(bitidx[3]), 
         .D(bitidx[0]), .Z(n38340)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(248[25:40])
    defparam i1_2_lut_rep_335_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_336_3_lut_4_lut (.A(cnt[0]), .B(cnt[1]), .C(n38402), 
         .D(cnt[5]), .Z(n38341)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_336_3_lut_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_adj_520 (.A(n486), .B(n6), .C(n1965), .D(n36406), 
         .Z(n36410)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_520.init = 16'hffec;
    LUT4 i1_4_lut_adj_521 (.A(bitidx[2]), .B(n3070), .C(n1963), .D(n3368), 
         .Z(n36406)) /* synthesis lut_function=(A (B+(C))+!A (C (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_521.init = 16'hf8a8;
    LUT4 i1_4_lut_adj_522 (.A(n5_adj_2258), .B(bitidx[3]), .C(n36392), 
         .D(n7), .Z(bitidx_3__N_195[3])) /* synthesis lut_function=(A+(B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_522.init = 16'heeea;
    LUT4 i1_4_lut_adj_523 (.A(n38359), .B(bitidx[3]), .C(n38401), .D(n38308), 
         .Z(n5_adj_2258)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_523.init = 16'h8882;
    LUT4 i1_3_lut_adj_524 (.A(n1965), .B(n36390), .C(n2895), .Z(n36392)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_3_lut_adj_524.init = 16'hecec;
    LUT4 i1_2_lut_rep_345_3_lut (.A(cnt[0]), .B(cnt[1]), .C(cnt[5]), .Z(n38350)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_345_3_lut.init = 16'hf7f7;
    LUT4 i23709_2_lut (.A(n68_adj_2233), .B(n32862), .Z(n2828)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23709_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_525 (.A(n38304), .B(n38302), .C(n3068), .D(n3070), 
         .Z(n36390)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_4_lut_adj_525.init = 16'hffec;
    LUT4 i25895_3_lut_4_lut (.A(cnt[0]), .B(cnt[1]), .C(cnt[5]), .D(cnt[6]), 
         .Z(n55)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam i25895_3_lut_4_lut.init = 16'hf008;
    LUT4 i23712_2_lut (.A(n71_adj_2234), .B(n32862), .Z(n2827)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23712_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_rep_397 (.A(cnt[4]), .B(cnt[2]), .C(cnt[3]), .Z(n38402)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_3_lut_rep_397.init = 16'h8080;
    LUT4 i1_2_lut_rep_341_4_lut (.A(cnt[4]), .B(cnt[2]), .C(cnt[3]), .D(n15), 
         .Z(n38346)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_rep_341_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_398 (.A(cnt[0]), .B(cnt[1]), .Z(n38403)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_rep_398.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_526 (.A(cnt[0]), .B(cnt[1]), .C(n15), .D(n103), 
         .Z(n13780)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_3_lut_4_lut_adj_526.init = 16'h0100;
    LUT4 i1_2_lut_rep_399 (.A(rx_ready), .B(n2352), .Z(n38404)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_rep_399.init = 16'h8888;
    LUT4 i1_4_lut_4_lut_4_lut (.A(rx_ready), .B(n2352), .C(n2355), .D(n38338), 
         .Z(fastclk_c_enable_14)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (D)+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_4_lut_4_lut.init = 16'hb8ff;
    LUT4 i1_3_lut_3_lut_adj_527 (.A(rx_ready), .B(n2352), .C(n2350), .Z(n10614)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_3_lut_3_lut_adj_527.init = 16'hd8d8;
    LUT4 i23026_2_lut_rep_400 (.A(n2353), .B(n2354), .Z(n38405)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23026_2_lut_rep_400.init = 16'heeee;
    LUT4 i31841_3_lut_4_lut (.A(n2353), .B(n2354), .C(n2352), .D(rx_ready), 
         .Z(n36546)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i31841_3_lut_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_401 (.A(n2354), .B(n2352), .Z(n38406)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_2_lut_rep_401.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_528 (.A(n2354), .B(n2352), .C(rx_ready), .D(reg_target[0]), 
         .Z(n13833)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_3_lut_4_lut_adj_528.init = 16'heee0;
    LUT4 i1_2_lut_rep_343_3_lut (.A(n2354), .B(n2352), .C(n2353), .Z(n38348)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_2_lut_rep_343_3_lut.init = 16'hfefe;
    LUT4 i23714_2_lut (.A(n74_adj_2235), .B(n32862), .Z(n2826)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23714_2_lut.init = 16'h2222;
    LUT4 i23717_2_lut (.A(n77_adj_2236), .B(n32862), .Z(n2825)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23717_2_lut.init = 16'h2222;
    LUT4 i23718_2_lut (.A(n80_adj_2237), .B(n32862), .Z(n2824)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23718_2_lut.init = 16'h2222;
    LUT4 i23721_2_lut (.A(n83_adj_2238), .B(n32862), .Z(n2823)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23721_2_lut.init = 16'h2222;
    LUT4 i23724_2_lut (.A(n86), .B(n32862), .Z(n2822)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23724_2_lut.init = 16'h2222;
    LUT4 i23727_2_lut (.A(n89), .B(n32862), .Z(n2821)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23727_2_lut.init = 16'h2222;
    LUT4 i23728_2_lut (.A(n92), .B(n32862), .Z(n2820)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23728_2_lut.init = 16'h2222;
    LUT4 i23731_2_lut (.A(n95), .B(n32862), .Z(n2819)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23731_2_lut.init = 16'h2222;
    LUT4 i23732_2_lut (.A(n98), .B(n32862), .Z(n2818)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23732_2_lut.init = 16'h2222;
    LUT4 i23745_2_lut (.A(n101), .B(n32862), .Z(n2817)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23745_2_lut.init = 16'h2222;
    LUT4 i23748_2_lut (.A(n104), .B(n32862), .Z(n2816)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23748_2_lut.init = 16'h2222;
    LUT4 i23751_2_lut (.A(n107), .B(n32862), .Z(n2815)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23751_2_lut.init = 16'h2222;
    LUT4 i23754_2_lut (.A(n110), .B(n32862), .Z(n2814)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23754_2_lut.init = 16'h2222;
    LUT4 i23757_2_lut (.A(n113), .B(n32862), .Z(n2813)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23757_2_lut.init = 16'h2222;
    LUT4 i23758_2_lut (.A(n116), .B(n32862), .Z(n2812)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23758_2_lut.init = 16'h2222;
    LUT4 i23767_2_lut (.A(n119), .B(n32862), .Z(n2811)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23767_2_lut.init = 16'h2222;
    LUT4 i23768_2_lut (.A(n122), .B(n32862), .Z(n2810)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23768_2_lut.init = 16'h2222;
    CCU2C add_26225_30 (.A0(gap[31]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n31205), 
          .S1(n1876));
    defparam add_26225_30.INIT0 = 16'h555f;
    defparam add_26225_30.INIT1 = 16'h0000;
    defparam add_26225_30.INJECT1_0 = "NO";
    defparam add_26225_30.INJECT1_1 = "NO";
    CCU2C add_26225_28 (.A0(gap[29]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[30]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31204), 
          .COUT(n31205));
    defparam add_26225_28.INIT0 = 16'h555f;
    defparam add_26225_28.INIT1 = 16'h555f;
    defparam add_26225_28.INJECT1_0 = "NO";
    defparam add_26225_28.INJECT1_1 = "NO";
    LUT4 tx_byte_0__bdd_3_lut_32992 (.A(tx_byte[0]), .B(tx_byte[1]), .C(bitidx[0]), 
         .Z(n37740)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;
    defparam tx_byte_0__bdd_3_lut_32992.init = 16'h3535;
    CCU2C add_26225_26 (.A0(gap[27]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[28]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31203), 
          .COUT(n31204));
    defparam add_26225_26.INIT0 = 16'h555f;
    defparam add_26225_26.INIT1 = 16'h555f;
    defparam add_26225_26.INJECT1_0 = "NO";
    defparam add_26225_26.INJECT1_1 = "NO";
    CCU2C add_26225_24 (.A0(gap[25]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[26]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31202), 
          .COUT(n31203));
    defparam add_26225_24.INIT0 = 16'h555f;
    defparam add_26225_24.INIT1 = 16'h555f;
    defparam add_26225_24.INJECT1_0 = "NO";
    defparam add_26225_24.INJECT1_1 = "NO";
    CCU2C add_26225_22 (.A0(gap[23]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[24]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31201), 
          .COUT(n31202));
    defparam add_26225_22.INIT0 = 16'h555f;
    defparam add_26225_22.INIT1 = 16'h555f;
    defparam add_26225_22.INJECT1_0 = "NO";
    defparam add_26225_22.INJECT1_1 = "NO";
    LUT4 i23769_2_lut (.A(n125), .B(n32862), .Z(n2809)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23769_2_lut.init = 16'h2222;
    pwm_led u_bar (.n5(n5), .fastclk_c(fastclk_c), .GND_net(GND_net), 
            .n39(n39_adj_2239), .distance({distance}), .VCC_net(VCC_net), 
            .n42(n42_adj_2240), .n83(n83), .n82(n82), .n81(n81), .n80(n80), 
            .n79(n79), .n78(n78), .n77(n77), .n76(n76), .n75(n75), 
            .n74(n74), .n73(n73), .n72(n72), .n71(n71), .n70(n70), 
            .n69(n69), .n68(n68), .n67(n67), .n66(n66), .n65(n65), 
            .n64(n64), .n63(n63), .n62(n62), .n61(n61), .n60(n60), 
            .n59(n59), .n58(n58), .n136(n136), .n51(n51_adj_2243), .n48(n48_adj_2242), 
            .n3556(n3556), .n75_adj_1(n75_adj_2251), .n45(n45_adj_2241), 
            .n66_adj_2(n66_adj_2216), .n63_adj_3(n63_adj_2218), .n60_adj_4(n60_adj_2246), 
            .n57(n57_adj_2245), .n72_adj_5(n72_adj_2217), .n69_adj_6(n69_adj_2222), 
            .n78_adj_7(n78_adj_2224), .n75_adj_8(n75_adj_2225), .n66_adj_9(n66_adj_2248), 
            .n63_adj_10(n63_adj_2247), .n84(n84_adj_2229), .n81_adj_11(n81_adj_2232), 
            .n90(n90), .n87(n87), .n96(n96), .n93(n93), .n102(n102), 
            .n99(n99), .n54(n54_adj_2244), .n69_adj_12(n69_adj_2249), 
            .n108(n108), .n105(n105), .n72_adj_13(n72_adj_2250), .n78_adj_14(n78_adj_2252), 
            .n114(n114), .n111(n111), .n81_adj_15(n81_adj_2253), .n120(n120), 
            .n117(n117), .n126(n126), .n123(n123), .n132(n132), .n129(n129), 
            .n138(n138), .n135(n135), .n141(n141), .led_c_3(led_c_3), 
            .led_c_2(led_c_2), .led_c_1(led_c_1), .led_c_0(led_c_0)) /* synthesis syn_module_defined=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(370[4] 375[3])
    CCU2C add_26225_20 (.A0(gap[21]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[22]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31200), 
          .COUT(n31201));
    defparam add_26225_20.INIT0 = 16'h555f;
    defparam add_26225_20.INIT1 = 16'h555f;
    defparam add_26225_20.INJECT1_0 = "NO";
    defparam add_26225_20.INJECT1_1 = "NO";
    CCU2C add_26225_18 (.A0(gap[19]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[20]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31199), 
          .COUT(n31200));
    defparam add_26225_18.INIT0 = 16'h555f;
    defparam add_26225_18.INIT1 = 16'h555f;
    defparam add_26225_18.INJECT1_0 = "NO";
    defparam add_26225_18.INJECT1_1 = "NO";
    CCU2C add_26225_16 (.A0(gap[17]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[18]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31198), 
          .COUT(n31199));
    defparam add_26225_16.INIT0 = 16'h555f;
    defparam add_26225_16.INIT1 = 16'h555f;
    defparam add_26225_16.INJECT1_0 = "NO";
    defparam add_26225_16.INJECT1_1 = "NO";
    LUT4 i23770_2_lut (.A(n128), .B(n32862), .Z(n2808)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23770_2_lut.init = 16'h2222;
    CCU2C add_26225_14 (.A0(gap[15]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[16]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31197), 
          .COUT(n31198));
    defparam add_26225_14.INIT0 = 16'h555f;
    defparam add_26225_14.INIT1 = 16'h555f;
    defparam add_26225_14.INJECT1_0 = "NO";
    defparam add_26225_14.INJECT1_1 = "NO";
    CCU2C add_26225_12 (.A0(gap[13]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[14]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31196), 
          .COUT(n31197));
    defparam add_26225_12.INIT0 = 16'h555f;
    defparam add_26225_12.INIT1 = 16'h555f;
    defparam add_26225_12.INJECT1_0 = "NO";
    defparam add_26225_12.INJECT1_1 = "NO";
    CCU2C add_26225_10 (.A0(gap[11]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[12]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31195), 
          .COUT(n31196));
    defparam add_26225_10.INIT0 = 16'h555f;
    defparam add_26225_10.INIT1 = 16'h555f;
    defparam add_26225_10.INJECT1_0 = "NO";
    defparam add_26225_10.INJECT1_1 = "NO";
    LUT4 i23771_2_lut (.A(n131), .B(n32862), .Z(n2807)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23771_2_lut.init = 16'h2222;
    CCU2C add_26225_8 (.A0(gap[9]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31194), 
          .COUT(n31195));
    defparam add_26225_8.INIT0 = 16'h555f;
    defparam add_26225_8.INIT1 = 16'h555f;
    defparam add_26225_8.INJECT1_0 = "NO";
    defparam add_26225_8.INJECT1_1 = "NO";
    CCU2C add_26225_6 (.A0(gap[7]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31193), 
          .COUT(n31194));
    defparam add_26225_6.INIT0 = 16'haaa0;
    defparam add_26225_6.INIT1 = 16'haaa0;
    defparam add_26225_6.INJECT1_0 = "NO";
    defparam add_26225_6.INJECT1_1 = "NO";
    CCU2C add_26225_4 (.A0(gap[5]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31192), 
          .COUT(n31193));
    defparam add_26225_4.INIT0 = 16'haaa0;
    defparam add_26225_4.INIT1 = 16'haaa0;
    defparam add_26225_4.INJECT1_0 = "NO";
    defparam add_26225_4.INJECT1_1 = "NO";
    LUT4 i23772_2_lut (.A(n134), .B(n32862), .Z(n2806)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23772_2_lut.init = 16'h2222;
    CCU2C add_26225_2 (.A0(gap[2]), .B0(gap[3]), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[4]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .COUT(n31192));
    defparam add_26225_2.INIT0 = 16'h000e;
    defparam add_26225_2.INIT1 = 16'haaa0;
    defparam add_26225_2.INJECT1_0 = "NO";
    defparam add_26225_2.INJECT1_1 = "NO";
    LUT4 i23773_2_lut (.A(n137), .B(n32862), .Z(n2805)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23773_2_lut.init = 16'h2222;
    LUT4 i23774_2_lut (.A(n140), .B(n32862), .Z(n2804)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23774_2_lut.init = 16'h2222;
    LUT4 i23775_2_lut (.A(n143), .B(n32862), .Z(n2803)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23775_2_lut.init = 16'h2222;
    LUT4 i23778_2_lut (.A(n146), .B(n32862), .Z(n2802)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23778_2_lut.init = 16'h2222;
    LUT4 i23779_2_lut (.A(n149), .B(n32862), .Z(n2801)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23779_2_lut.init = 16'h2222;
    LUT4 i23784_2_lut (.A(n152), .B(n32862), .Z(n2800)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23784_2_lut.init = 16'h2222;
    LUT4 i23785_2_lut (.A(n155), .B(n32862), .Z(n2799)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23785_2_lut.init = 16'h2222;
    LUT4 i23786_2_lut (.A(n158), .B(n32862), .Z(n2798)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23786_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_529 (.A(reg_target[4]), .B(rx_ready), .C(n34245), 
         .D(n38405), .Z(reg_target_7__N_247[4])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_529.init = 16'heca0;
    LUT4 i1_4_lut_adj_530 (.A(n2960), .B(rx_ready), .C(n38405), .D(n2352), 
         .Z(n34245)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(38[9:17])
    defparam i1_4_lut_adj_530.init = 16'hfbfa;
    LUT4 i1_4_lut_adj_531 (.A(reg_target[3]), .B(rx_ready), .C(n34248), 
         .D(n13), .Z(reg_target_7__N_247[3])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_4_lut_adj_531.init = 16'heca0;
    LUT4 i1_4_lut_adj_532 (.A(n2960), .B(rx_ready), .C(n2352), .D(n38405), 
         .Z(n34248)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_4_lut_adj_532.init = 16'hfbfa;
    LUT4 i1_4_lut_adj_533 (.A(rx_ready), .B(reg_target[2]), .C(n38342), 
         .D(n38339), .Z(reg_target_7__N_247[2])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_4_lut_adj_533.init = 16'heca0;
    LUT4 i1_4_lut_adj_534 (.A(reg_target[1]), .B(n38348), .C(n2960), .D(rx_ready), 
         .Z(reg_target_7__N_247[1])) /* synthesis lut_function=(A (B+(C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(304[13] 360[20])
    defparam i1_4_lut_adj_534.init = 16'heca8;
    LUT4 i23601_2_lut (.A(reg_target[7]), .B(n27539), .Z(n2748)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23601_2_lut.init = 16'h8888;
    CCU2C add_26226_10 (.A0(gap[9]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[10]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30551), 
          .COUT(n30552));
    defparam add_26226_10.INIT0 = 16'h555f;
    defparam add_26226_10.INIT1 = 16'h555f;
    defparam add_26226_10.INJECT1_0 = "NO";
    defparam add_26226_10.INJECT1_1 = "NO";
    LUT4 i23598_2_lut (.A(reg_target[3]), .B(n27539), .Z(n2744)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i23598_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_535 (.A(n27539), .B(reg_target[2]), .Z(n2743)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_535.init = 16'h8888;
    LUT4 i1_2_lut_adj_536 (.A(n36), .B(n34), .Z(cnt_15__N_167[15])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_536.init = 16'h8888;
    LUT4 i1_2_lut_adj_537 (.A(n39), .B(n34), .Z(cnt_15__N_167[14])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_537.init = 16'h8888;
    LUT4 i1_2_lut_adj_538 (.A(n42), .B(n34), .Z(cnt_15__N_167[13])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_538.init = 16'h8888;
    LUT4 i1_2_lut_adj_539 (.A(n45), .B(n34), .Z(cnt_15__N_167[12])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_539.init = 16'h8888;
    LUT4 i1_2_lut_adj_540 (.A(n48), .B(n34), .Z(cnt_15__N_167[11])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_540.init = 16'h8888;
    LUT4 i1_2_lut_adj_541 (.A(n51), .B(n34), .Z(cnt_15__N_167[10])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_541.init = 16'h8888;
    LUT4 i1_2_lut_adj_542 (.A(n54), .B(n34), .Z(cnt_15__N_167[9])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_542.init = 16'h8888;
    LUT4 i1_2_lut_adj_543 (.A(n57), .B(n34), .Z(cnt_15__N_167[8])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_543.init = 16'h8888;
    LUT4 i1_2_lut_adj_544 (.A(n60_adj_2226), .B(n34), .Z(cnt_15__N_167[7])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_544.init = 16'h8888;
    LUT4 i1_2_lut_adj_545 (.A(n63_adj_2223), .B(n34), .Z(cnt_15__N_167[6])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_545.init = 16'h8888;
    CCU2C _add_1_1298_add_4_17 (.A0(distance[15]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30497), .S0(n5));
    defparam _add_1_1298_add_4_17.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_17.INIT1 = 16'h0000;
    defparam _add_1_1298_add_4_17.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_546 (.A(n66_adj_2230), .B(n34), .Z(cnt_15__N_167[5])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_546.init = 16'h8888;
    LUT4 i1_2_lut_adj_547 (.A(n69_adj_2228), .B(n34), .Z(cnt_15__N_167[4])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_547.init = 16'h8888;
    LUT4 i1_2_lut_adj_548 (.A(n72_adj_2227), .B(n34), .Z(cnt_15__N_167[3])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_548.init = 16'h8888;
    LUT4 i1_2_lut_adj_549 (.A(n75_adj_2219), .B(n34), .Z(cnt_15__N_167[2])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_549.init = 16'h8888;
    LUT4 i1_2_lut_adj_550 (.A(n78_adj_2220), .B(n34), .Z(cnt_15__N_167[1])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i1_2_lut_adj_550.init = 16'h8888;
    LUT4 i6640_4_lut (.A(n1969), .B(n1959), .C(n38304), .D(n33465), 
         .Z(n10580)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(116[13] 301[20])
    defparam i6640_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_551 (.A(n36608), .B(n36664), .C(n36614), .D(n36596), 
         .Z(n34576)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_adj_551.init = 16'hfffb;
    LUT4 i1_4_lut_adj_552 (.A(msb[7]), .B(lsb[6]), .C(msb[3]), .D(lsb[7]), 
         .Z(n36608)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_adj_552.init = 16'hfffe;
    LUT4 i31831_2_lut (.A(lsb[2]), .B(lsb[4]), .Z(n36664)) /* synthesis lut_function=(A (B)) */ ;
    defparam i31831_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_553 (.A(lsb[3]), .B(n36610), .C(n36600), .D(msb[5]), 
         .Z(n36614)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_adj_553.init = 16'hfffe;
    LUT4 i1_2_lut_adj_554 (.A(lsb[1]), .B(msb[2]), .Z(n36596)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_adj_554.init = 16'heeee;
    LUT4 i1_4_lut_adj_555 (.A(lsb[0]), .B(msb[4]), .C(lsb[5]), .D(msb[0]), 
         .Z(n36610)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_4_lut_adj_555.init = 16'hfffe;
    LUT4 i1_2_lut_adj_556 (.A(msb[1]), .B(msb[6]), .Z(n36600)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_adj_556.init = 16'heeee;
    LUT4 i1_2_lut_adj_557 (.A(rx_ready), .B(n2350), .Z(n36620)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(82[12] 362[8])
    defparam i1_2_lut_adj_557.init = 16'h8888;
    LUT4 n1965_bdd_4_lut_32765 (.A(n1965), .B(n38327), .C(n38347), .D(n1964), 
         .Z(n27539)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam n1965_bdd_4_lut_32765.init = 16'h0002;
    PFUMX i22364 (.BLUT(n28), .ALUT(n26314), .C0(n1960), .Z(rx_remaining_1__N_292[0]));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    VLO i1 (.Z(GND_net));
    PFUMX i32483 (.BLUT(n38122), .ALUT(n38121), .C0(n38358), .Z(n38123));
    PFUMX i32481 (.BLUT(n38117), .ALUT(n38116), .C0(n1967), .Z(n38118));
    PFUMX i32514 (.BLUT(n38428), .ALUT(n38429), .C0(bitidx[2]), .Z(n38430));
    PFUMX i32512 (.BLUT(n38425), .ALUT(n38426), .C0(n1965), .Z(n38427));
    CCU2C add_26226_8 (.A0(gap[7]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[8]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30550), 
          .COUT(n30551));
    defparam add_26226_8.INIT0 = 16'h555f;
    defparam add_26226_8.INIT1 = 16'h555f;
    defparam add_26226_8.INJECT1_0 = "NO";
    defparam add_26226_8.INJECT1_1 = "NO";
    CCU2C _add_1_1298_add_4_15 (.A0(distance[14]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[15]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30496), .COUT(n30497), .S0(n42_adj_2240), 
          .S1(n39_adj_2239));
    defparam _add_1_1298_add_4_15.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_15.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_15.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_15.INJECT1_1 = "NO";
    PFUMX i32510 (.BLUT(n38422), .ALUT(n38423), .C0(n38324), .Z(n32862));
    PFUMX i32508 (.BLUT(n38419), .ALUT(n38420), .C0(bitidx[0]), .Z(n38421));
    CCU2C _add_1_1298_add_4_13 (.A0(distance[12]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[13]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30495), .COUT(n30496), .S0(n48_adj_2242), 
          .S1(n45_adj_2241));
    defparam _add_1_1298_add_4_13.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_13.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_13.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_13.INJECT1_1 = "NO";
    CCU2C _add_1_1298_add_4_11 (.A0(distance[10]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[11]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30494), .COUT(n30495), .S0(n54_adj_2244), 
          .S1(n51_adj_2243));
    defparam _add_1_1298_add_4_11.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_11.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_11.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_11.INJECT1_1 = "NO";
    CCU2C add_26226_6 (.A0(gap[5]), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(gap[6]), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30549), 
          .COUT(n30550));
    defparam add_26226_6.INIT0 = 16'h555f;
    defparam add_26226_6.INIT1 = 16'h555f;
    defparam add_26226_6.INJECT1_0 = "NO";
    defparam add_26226_6.INJECT1_1 = "NO";
    CCU2C _add_1_1298_add_4_9 (.A0(distance[8]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[9]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n30493), .COUT(n30494), .S0(n60_adj_2246), 
          .S1(n57_adj_2245));
    defparam _add_1_1298_add_4_9.INIT0 = 16'h555f;
    defparam _add_1_1298_add_4_9.INIT1 = 16'h555f;
    defparam _add_1_1298_add_4_9.INJECT1_0 = "NO";
    defparam _add_1_1298_add_4_9.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module pwm_led
//

module pwm_led (n5, fastclk_c, GND_net, n39, distance, VCC_net, 
            n42, n83, n82, n81, n80, n79, n78, n77, n76, n75, 
            n74, n73, n72, n71, n70, n69, n68, n67, n66, n65, 
            n64, n63, n62, n61, n60, n59, n58, n136, n51, 
            n48, n3556, n75_adj_1, n45, n66_adj_2, n63_adj_3, n60_adj_4, 
            n57, n72_adj_5, n69_adj_6, n78_adj_7, n75_adj_8, n66_adj_9, 
            n63_adj_10, n84, n81_adj_11, n90, n87, n96, n93, n102, 
            n99, n54, n69_adj_12, n108, n105, n72_adj_13, n78_adj_14, 
            n114, n111, n81_adj_15, n120, n117, n126, n123, n132, 
            n129, n138, n135, n141, led_c_3, led_c_2, led_c_1, 
            led_c_0) /* synthesis syn_module_defined=1 */ ;
    input n5;
    input fastclk_c;
    input GND_net;
    input n39;
    input [15:0]distance;
    input VCC_net;
    input n42;
    output n83;
    output n82;
    output n81;
    output n80;
    output n79;
    output n78;
    output n77;
    output n76;
    output n75;
    output n74;
    output n73;
    output n72;
    output n71;
    output n70;
    output n69;
    output n68;
    output n67;
    output n66;
    output n65;
    output n64;
    output n63;
    output n62;
    output n61;
    output n60;
    output n59;
    output n58;
    output n136;
    input n51;
    input n48;
    input n3556;
    input n75_adj_1;
    input n45;
    input n66_adj_2;
    input n63_adj_3;
    input n60_adj_4;
    input n57;
    input n72_adj_5;
    input n69_adj_6;
    input n78_adj_7;
    input n75_adj_8;
    input n66_adj_9;
    input n63_adj_10;
    input n84;
    input n81_adj_11;
    input n90;
    input n87;
    input n96;
    input n93;
    input n102;
    input n99;
    input n54;
    input n69_adj_12;
    input n108;
    input n105;
    input n72_adj_13;
    input n78_adj_14;
    input n114;
    input n111;
    input n81_adj_15;
    input n120;
    input n117;
    input n126;
    input n123;
    input n132;
    input n129;
    input n138;
    input n135;
    input n141;
    output led_c_3;
    output led_c_2;
    output led_c_1;
    output led_c_0;
    
    wire fastclk_c /* synthesis SET_AS_NETWORK=fastclk_c, is_clock=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/top.v(6[16:23])
    
    wire n1744;
    wire [31:0]n1808;
    
    wire n38295, n1846, n35744, n30608, n13631, n28090, n1748, 
        n1747;
    wire [31:0]n1907;
    
    wire n30609, n30810, n13547, n28588;
    wire [31:0]n3194;
    
    wire n3135, n3134;
    wire [31:0]n3293;
    
    wire n30811, n38331;
    wire [31:0]n1709;
    wire [31:0]n2;
    
    wire n1746, n28568, n13550;
    wire [31:0]n2897;
    
    wire n2832, n2931;
    wire [31:0]n1709_adj_2160;
    wire [31:0]n35;
    
    wire n1744_adj_520, n2848, n2947, n30607, n1750, n1749, n30606, 
        n1752, n1751, n30688, n13590, n28440;
    wire [31:0]n2204;
    
    wire n38275, n38274;
    wire [31:0]n2303;
    wire [14:0]pwm_cnt;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(27[19:26])
    
    wire n14116;
    wire [14:0]n50;
    
    wire n2838, n2937, n28434, n13620;
    wire [31:0]n3293_adj_2161;
    
    wire n3241, n3340, n30547, n13629, n28492, n3227;
    wire [31:0]n3392;
    
    wire n3246, n3345, n30546, n38190, n3228, n30605, n1754, n1753;
    wire [10:0]n3568;
    
    wire n3549;
    wire [10:0]n36;
    
    wire n30604, n12154, n38307, n30687, n2141, n2140;
    wire [31:0]duty0_14__N_426;
    
    wire n594, n30809, n3137, n3136, n2853;
    wire [31:0]n2897_adj_2162;
    
    wire n38226, n2951, n34692, n3233, n3332, n30808, n3139, n3138, 
        n2842, n2940, n35208, n3547, n3548, n587, n28307, n13598, 
        n27382, n3, n2834, n38220, n38224, n3550, n38225, n3546, 
        n30545, n3231, n3230;
    wire [14:0]duty0;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    
    wire n12416;
    wire [14:0]duty0_14__N_410;
    
    wire n3454, n3551, n38179, n3449, n3458, n38175, n30544, n3233_adj_522, 
        n3232, n34756, n33580, n34758, n39_adj_523, n38229, n2930;
    wire [14:0]duty1;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[26:31])
    wire [14:0]duty1_14__N_458;
    wire [14:0]duty2;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[33:38])
    wire [14:0]duty2_14__N_473;
    wire [14:0]duty3;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[40:45])
    wire [14:0]duty3_14__N_488;
    
    wire n30603;
    wire [31:0]n1412;
    
    wire n30686, n2143, n2142, n30543, n3235, n3234, n30602, n3435, 
        n34752, n34740, n3437, n2838_adj_525, n2937_adj_526, n586, 
        n2843, n2942, n3446, n31, n34746, n3434, n30807, n3141, 
        n3140, n30806, n38201, n3142, n30979, n13624, n28462;
    wire [31:0]n2699;
    
    wire n2643, n2642;
    wire [31:0]n2798;
    
    wire n30980;
    wire [31:0]n4540;
    
    wire n31386, n3443, n3440, n3436, n3441, n344, n30978, n2645, 
        n2644, n38238, n2939, n334, n2847, n2946, n338, n30977, 
        n2647, n2646, n3351;
    wire [31:0]n3392_adj_2163;
    
    wire n3359, n3450, n30976, n2649, n2648, n30601, n345, n30685, 
        n38277, n2144, n2839, n2938, n30805, n3145, n3144, n30804, 
        n3147, n3146, n30975, n2651, n2650, n585, n341, n3353, 
        n3452, n30684, n2147, n2146, n30542, n3237, n3236, n30541, 
        n3239, n3238, n2841, n30600, n30540, n3241_adj_532, n3240, 
        n30539, n3243, n3242, n2854, n2953, n3354, n3453, n2835, 
        n2934, n2832_adj_534, n2931_adj_535, n30599, n30683, n2149, 
        n2148, n38187, n3451, n37665, n37664, n38177, n37666, 
        n30597, n13600, n28359, n1842, n1841;
    wire [31:0]n2006;
    
    wire n3334, n3433, n3250, n3349, n38191, n3330, n2836, n2935, 
        n3235_adj_539, n30538, n3245, n3244, n3347, n2845, n2944, 
        n3346, n3438, n3339, n2844, n2943, n3237_adj_542, n3336, 
        n3335, n30596, n38291, n38290, n30682, n2151, n2150, n30803, 
        n3149, n3148, n3338, n30595, n1845, n38235, n2936, n3344, 
        n2833, n2932, n30537, n3247, n3246_adj_548, n3244_adj_551, 
        n3343, n30594, n1848, n1847, n30681, n2153, n38278, n30536, 
        n3249, n3248, n30593, n1850, n1849, n30592, n38292, n1851, 
        n30680, n337, n2154, n30802, n38202, n3150, n30974, n2653, 
        n2652, n30535, n38196, n3250_adj_554, n2846, n2945, n593, 
        n2954, n3341, n3337, n3342, n38237, n30973, n342, n2654, 
        n3447, n30534, n3253, n3252, n3240_adj_561, n34976, n38059, 
        n3428, n3444, n38186, n3425, n28528, n13610;
    wire [31:0]n3293_adj_2164;
    
    wire n3240_adj_564, n3339_adj_565, n38184, n3236_adj_568, n2848_adj_570, 
        n2947_adj_571, n30533, n348, n3254, n3326, n2849, n2948, 
        n38163, n1;
    wire [32:0]n197;
    
    wire n2983, n13790;
    wire [32:0]n89;
    
    wire n30801, n3153, n3152, n3348, n3229, n3328, n2850, n2949, 
        n3243_adj_580, n38178, n2851, n2950, n36114, n36120, n36110, 
        n36116, n36112, n36090, n35824, n35786, n28176, n3545, 
        n598, n3228_adj_582, n3327, n2039, n34486, n36046, n2042, 
        n13605, n3227_adj_584, n2045, n2043, n2044, n2041, n38232, 
        n38228, n2845_adj_585, n35452, n30800, n347, n3154, n343, 
        n30679, n28263;
    wire [31:0]n2105;
    
    wire n28468, n13622, n2047, n28247, n2048, n2049, n30971, 
        n13625, n28456;
    wire [31:0]n2600;
    
    wire n2535, n2534, n38198, n30970, n2537, n2536, n2051, n2050, 
        n27986, n2052, n38227, n336, n2053, n2054, n3242_adj_588, 
        n2739, n38222, n30969, n2539, n2538, n16_adj_589, n22, 
        n36923, n24, n30591, n1854, n1853, n30528;
    wire [31:0]n38;
    
    wire n2754, n2853_adj_591, n30968, n2541, n2540, n2741, n2840, 
        n2733, n2832_adj_592, n30678, n2040, n30677, n30590, n583, 
        n30967, n2543, n2542, n30799, n13548, n28578;
    wire [31:0]n3095;
    
    wire n3029, n30798, n38211, n38212, n35684, n35678, n2545, 
        n35680, n30527, n2544, n2746, n3254_adj_597, n30797, n3033, 
        n3032, n30796, n3035, n3034, n2546, n3247_adj_599, n38316, 
        n2854_adj_601, n30676, n30966, n38317, n30795, n3037, n3036, 
        n2548, n28299, n2547, n2549, n3242_adj_603, n3341_adj_604, 
        n2551, n2550, n28048, n2552, n30794, n3039, n3038, n341_adj_605, 
        n2553, n2554, n30965, n3251, n3350, n16_adj_607, n22_adj_608, 
        n36866, n24_adj_609, n2748, n2847_adj_610, n2734, n38219, 
        n30675, n38281, n3231_adj_612, n3330_adj_613, n597, n2732, 
        n2831, n2747, n2846_adj_615, n30964, n30963, n30674, n30962, 
        n30961, n30793, n3041, n3040, n2742, n2841_adj_616, n3248_adj_618, 
        n2753, n2852, n30960, n13627, n28446;
    wire [31:0]n2501;
    
    wire n38254, n2736, n2835_adj_619, n2743, n2842_adj_620, n3249_adj_622, 
        n30792, n3043, n3042, n3239_adj_624, n30959, n2437, n2436, 
        n16_adj_625, n22_adj_626, n36809, n24_adj_627, n30673, n30791, 
        n3045, n3044, n2737, n2836_adj_628, n3234_adj_630, n3333, 
        n2750, n2849_adj_631, n3327_adj_632, n3332_adj_633, n3345_adj_634, 
        n3335_adj_635, n37516, n2751, n2850_adj_636, n2744, n2843_adj_637, 
        n3238_adj_639, n38398, n38397, n38396, n36909, n36010, n36000;
    wire [14:0]n4990;
    
    wire n36008, n35982, n3046, n35992, n36002, n2735, n2834_adj_640, 
        n3245_adj_642, n38233, n2839_adj_643, n2738, n2837, n3047, 
        n28496, n3048, n3049, n28522, n13614, n38189, n3051, n3050, 
        n28190, n3052, n30526, n346, n3053, n3054, n2749, n2848_adj_646, 
        n2752, n2851_adj_647, n2732_adj_648;
    wire [31:0]n2798_adj_2165;
    
    wire n38239, n35428, n2734_adj_650;
    wire [31:0]n2798_adj_2166;
    
    wire n38240, n36188, n16_adj_652, n22_adj_653, n36752, n24_adj_654;
    wire [31:0]n3194_adj_2167;
    
    wire n3154_adj_656, n3253_adj_657, n30525, n3138_adj_661, n3237_adj_662, 
        n2736_adj_663, n2839_adj_665, n36196, n347_adj_667, n3254_adj_668, 
        n38234, n35376, n30672, n592, n3152_adj_671, n3251_adj_672, 
        n3137_adj_674, n3236_adj_675, n343_adj_677, n38322, n3131, 
        n38182, n30671, n2641, n35384, n30589, n13604, n28333, 
        n1940;
    wire [31:0]n2105_adj_2168;
    
    wire n38192, n3228_adj_682, n3142_adj_684, n3241_adj_685, n3135_adj_687, 
        n3234_adj_688, n30958, n2439, n2438, n30790, n30789, n30788, 
        n30957, n2441, n38255, n30669, n38306, n30787, n3144_adj_691, 
        n3243_adj_692, n2635, n3149_adj_694, n3248_adj_695, n30786, 
        n30956, n2443, n2442, n3150_adj_697, n3249_adj_698, n30955, 
        n2445, n2444, n30588, n1942, n1941, n30524, n30954, n2447, 
        n2446, n3151, n3250_adj_704, n30668, n30953, n2449, n2448, 
        n30952, n2451, n2450, n38241, n30784, n13549, n28574;
    wire [31:0]n2996;
    
    wire n2930_adj_706, n30667, n30587, n1944, n1943, n30783, n38221, 
        n2932_adj_709, n30782, n2935_adj_710, n2934_adj_711, n30666, 
        n2638, n30951, n2453, n2452, n30586, n1946, n1945, n30523, 
        n3153_adj_717, n3252_adj_718, n3245_adj_720, n3344_adj_721, 
        n38193, n3229_adj_723, n28562, n13640;
    wire [31:0]n1709_adj_2169;
    
    wire n331, n1753_adj_724, n2636, n30950, n340, n2454, n3128, 
        n3227_adj_726, n30585, n1948, n1947, n3141_adj_730, n30948, 
        n13630, n28442;
    wire [31:0]n2402;
    
    wire n2337, n2336, n30665, n30584, n1950, n1949, n3143, n2639, 
        n30664, n3246_adj_736, n38392, n38391, n38390, n36852, n2634, 
        n30781, n2936_adj_737, n2640, n30583, n1952, n1951, n30947, 
        n2339, n2338, n35556, n35540, n30780, n2939_adj_740, n2938_adj_741, 
        n30779, n2941, n2940_adj_742, n35552, n35538, n30582, n1954, 
        n1953, n28309, n28052, n30778, n2943_adj_745, n2942_adj_746, 
        n30946, n2341, n2340, n30777, n2945_adj_747, n2944_adj_748, 
        n30663, n30945, n38262, n2342, n30522, n38194, n30944, 
        n2345, n2344, n2637, n3139_adj_753, n3238_adj_754, n30661, 
        n13613, n28526;
    wire [31:0]n2006_adj_2170;
    
    wire n1941_adj_756, n1940_adj_758, n30776, n2946_adj_759, n2738_adj_760, 
        n35424, n2742_adj_762, n2842_adj_764, n36186, n28512, n13602, 
        n3133, n3232_adj_766, n3146_adj_768, n3147_adj_770, n3140_adj_772, 
        n3239_adj_773, n2753_adj_774, n34684, n30943, n2347, n2346, 
        n30660, n1943_adj_777, n1942_adj_779, n2741_adj_780, n35434, 
        n30659, n1945_adj_783, n1944_adj_785, n37667, n28373, n13626, 
        n38386, n38385, n38384, n36795, n30775, n2949_adj_786, n2948_adj_787, 
        n30521, n3136_adj_791, n3235_adj_792, n3134_adj_794, n3233_adj_795, 
        n2745, n2737_adj_798, n30658, n1947_adj_800, n1946_adj_802, 
        n30581, n584, n3145_adj_806, n3244_adj_807, n3336_adj_808, 
        n43, n30942, n2349, n2348, n3148_adj_810, n3247_adj_811, 
        n30941, n2351, n2350, n30940, n2353, n2352, n30939, n339, 
        n2354, n3330_adj_812, n55, n38380, n38379, n38378, n36738, 
        n2735_adj_814, n2739_adj_816, n35742, n2746_adj_818, n28174, 
        n27898, n30774, n2951_adj_819, n2950_adj_820, n36154, n36144, 
        n36148, n36134, n36146, n2744_adj_822, n3130, n38197, n2747_adj_824, 
        n38242, n30657, n1949_adj_827, n1948_adj_829, n30773, n2953_adj_830, 
        n2952, n333, n28502, n28202, n30656, n1951_adj_833, n1950_adj_835, 
        n30772, n2954_adj_836, n30655, n1953_adj_838, n1952_adj_840, 
        n35624, n12_adj_841, n26_adj_842, n36947, n28, n30938, n13633, 
        n28430;
    wire [31:0]n2303_adj_2171;
    
    wire n2237, n38305, n38321, n30579, n13595, n28407, n2040_adj_844, 
        n2039_adj_845;
    wire [31:0]n2204_adj_2172;
    
    wire n30578, n2042_adj_849, n2041_adj_850, n35620, n35608, n38332, 
        n30937, n2239, n2238, n30771, n2831_adj_857, n30936, n2241, 
        n2240, n2740, n28315, n30654, n335, n1954_adj_863, n30935, 
        n2243, n2242, n28058, n36338, n28249, n30520, n27990, 
        n30770, n38230, n38333, n38244, n30934, n2245, n2244, 
        n36927, n30653, n38289, n28321;
    wire [31:0]n1907_adj_2173;
    
    wire n1841_adj_874, n3339_adj_875, n37, n30933, n2247, n2246, 
        n30769, n38231, n2834_adj_880, n30932, n2249, n2248, n2733_adj_884, 
        n30768, n2837_adj_886, n2836_adj_888, n2743_adj_890, n38374, 
        n38376, n36891, n2742_adj_892, n38334, n30767, n30931, n2251, 
        n2250, n30766, n38236, n2840_adj_899, n30930, n2253, n2252, 
        n30765, n2843_adj_903, n30577, n2044_adj_905, n38280, n35516, 
        n35514, n30519, n2748_adj_911, n28317, n30929, n338_adj_913, 
        n2254, n28060, n38335, n30764, n2845_adj_917, n2844_adj_919, 
        n30518, n35694, n35692, n2045_adj_922, n2046, n2047_adj_923, 
        n28168, n2048_adj_924, n2049_adj_925, n2051_adj_926, n2050_adj_927, 
        n27890, n2052_adj_928, n30927, n13634, n28412;
    wire [31:0]n2204_adj_2174;
    
    wire n2139, n2138, n2053_adj_931, n2054_adj_932, n30763, n2847_adj_934, 
        n2846_adj_936, n3132;
    wire [31:0]n3194_adj_2175;
    
    wire n38199, n35264, n36208, n36202, n30762, n2849_adj_939, 
        n2749_adj_941, n2750_adj_943, n2754_adj_945, n36204, n38246, 
        n3030;
    wire [31:0]n3095_adj_2176;
    
    wire n38195, n35342, n28508, n2751_adj_950, n2851_adj_951, n2850_adj_952, 
        n28210, n2852_adj_953, n2853_adj_954, n2854_adj_955, n28554, 
        n13551, n1844, n1846_adj_956, n1842_adj_957, n36346, n1847_adj_958, 
        n28257, n1848_adj_959, n1849_adj_960, n30652, n1843, n1851_adj_963, 
        n1850_adj_964, n28006, n1852, n2743_adj_966, n1853_adj_967, 
        n1854_adj_968, n30576, n30575, n30651, n1845_adj_974, n30517, 
        n30516, n35660, n35658, n2141_adj_983, n2143_adj_984, n2146_adj_985, 
        n2144_adj_986, n30515, n2751_adj_989, n2142_adj_990, n2145, 
        n2140_adj_991, n2148_adj_992, n28329, n2147_adj_993, n2149_adj_994, 
        n2151_adj_995, n2150_adj_996, n28070, n2152, n2735_adj_998, 
        n30761, n337_adj_1001, n2153_adj_1002, n2154_adj_1003, n30574, 
        n30926, n30650, n30925, n30760, n36160, n36178, n36176, 
        n30573, n30924, n2737_adj_1018, n36174, n36168, n2733_adj_1019, 
        n30759, n30572, n30571, n30649, n30648, n33356, n38164, 
        n60_adj_1030, n2744_adj_1032, n2745_adj_1033, n2746_adj_1034, 
        n2739_adj_1035, n2741_adj_1036, n2754_adj_1038, n2747_adj_1039, 
        n28510, n2748_adj_1040, n2749_adj_1041, n2753_adj_1043, n3031, 
        n35338, n2750_adj_1046, n28214, n2752_adj_1047, n2045_adj_1048, 
        n35716, n35714, n2043_adj_1049, n13635, n2044_adj_1050, n2040_adj_1051, 
        n2046_adj_1052, n2042_adj_1053, n3033_adj_1055, n35348, n2048_adj_1058, 
        n28337, n2047_adj_1059, n2049_adj_1060, n28401, n2051_adj_1061, 
        n2050_adj_1062, n27972, n2052_adj_1063, n336_adj_1064, n2053_adj_1065, 
        n2054_adj_1066, n35960, n13653, n35834, n1750_adj_1073, n34329, 
        n28287, n35830, n1754_adj_1076, n30647, n36870, n28518, 
        n13617, n38245, n30757, n38243, n30756, n30755, n30646, 
        n30754, n2738_adj_1089, n30923;
    wire [31:0]n3392_adj_2177;
    
    wire n37486, n38370, n38372, n36834, n36943, n30922, n30921, 
        n30920, n30919, n30918;
    wire [31:0]n2105_adj_2178;
    
    wire n38273, n30917, n2041_adj_1109, n30753, n3347_adj_1112, n21_adj_1113, 
        n3341_adj_1114, n33, n3040_adj_1116, n30916, n35706, n1945_adj_1119, 
        n1940_adj_1120, n1942_adj_1121, n13636, n30915, n1944_adj_1125, 
        n1941_adj_1126, n1943_adj_1127, n1946_adj_1128, n38249, n35074, 
        n30914, n1948_adj_1132, n28343, n1947_adj_1133, n1949_adj_1134, 
        n28389, n30644;
    wire [31:0]n1808_adj_2179;
    
    wire n1743, n1742, n30643, n1745, n346_adj_1140, n30752, n30913, 
        n1951_adj_1143, n1950_adj_1144, n28080, n1952_adj_1145, n2635_adj_1146;
    wire [31:0]n2699_adj_2180;
    
    wire n38248, n35410, n30912, n335_adj_1150, n1953_adj_1151, n1954_adj_1152, 
        n30751, n36232, n36226, n2635_adj_1153, n2636_adj_1154, n13552, 
        n2633;
    wire [31:0]n2699_adj_2181;
    
    wire n38247, n2641_adj_1156, n36228, n36220, n2646_adj_1157, n30911, 
        n30750, n30910, n30749, n2640_adj_1162, n2634_adj_1163, n2639_adj_1164, 
        n2638_adj_1165, n30748, n2637_adj_1166, n2643_adj_1167, n2644_adj_1168, 
        n2647_adj_1169, n28514, n2648_adj_1170, n2649_adj_1171, n28544, 
        n2651_adj_1172, n2650_adj_1173, n28218, n2652_adj_1174, n3036_adj_1176, 
        n12_adj_1177, n26_adj_1178, n28_adj_1179, n3050_adj_1181, n3053_adj_1183, 
        n342_adj_1184, n2653_adj_1185, n2654_adj_1186, n1841_adj_1187, 
        n1844_adj_1188, n1843_adj_1189, n1842_adj_1190, n35726, n1848_adj_1191, 
        n28351, n1847_adj_1192, n1849_adj_1193, n28377, n1851_adj_1194, 
        n1850_adj_1195, n28086, n1852_adj_1196, n30908;
    wire [31:0]n2006_adj_2182;
    
    wire n334_adj_1199, n1853_adj_1200, n1854_adj_1201, n2637_adj_1202, 
        n35402, n36813, n30642, n1747_adj_1206, n1746_adj_1208, n30747, 
        n3343_adj_1209, n3347_adj_1210, n37505, n30746, n30641, n1749_adj_1212, 
        n38297, n2653_adj_1214, n34654, n3045_adj_1217, n30907, n30906, 
        n30905, n30745, n30744, n3038_adj_1227, n38366, n38368, 
        n36777, n36939, n30640, n1751_adj_1229, n30904, n36308, 
        n36302, n2545_adj_1233, n2546_adj_1234, n13553, n2539_adj_1235, 
        n36304, n2537_adj_1236, n2536_adj_1237, n2540_adj_1238, n2544_adj_1239, 
        n2541_adj_1240, n2542_adj_1241, n30903, n2538_adj_1245, n2535_adj_1246, 
        n2543_adj_1247, n2534_adj_1248, n2547_adj_1249, n28226, n2548_adj_1250, 
        n2549_adj_1251, n28331, n30743, n30902, n30742, n2551_adj_1259, 
        n2550_adj_1260, n27956, n2552_adj_1261, n30901, n3054_adj_1265, 
        n30741, n30639, n1753_adj_1268, n1752_adj_1270, n30900, n38283;
    wire [31:0]n1907_adj_2183;
    
    wire n2553_adj_1272, n2554_adj_1273, n3346_adj_1276, n23_adj_1277;
    wire [31:0]n1610;
    
    wire n33572, n34842, n34848, n34838, n34816, n34846, n30899, 
        n38282, n28281, n13628;
    wire [31:0]n3095_adj_2184;
    
    wire n38216, n3151_adj_1294, n3044_adj_1296, n3143_adj_1297, n34732, 
        n34782, n1650, n28104, n1647, n1648, n1649, n332, n1653, 
        n1654, n330, n28558, n329, n1652, n1350, n1351, n1352, 
        n1353, n1448, n1646, n3042_adj_1299, n2642_adj_1302, n3326_adj_1304, 
        n63_adj_1305, n36756, n3328_adj_1306, n38173, n3338_adj_1307, 
        n37487, n38362, n38364, n36720, n36935, n36286, n2437_adj_1310, 
        n36270, n2445_adj_1311, n13554, n2438_adj_1312, n36282, n36268, 
        n2446_adj_1313, n3029_adj_1316, n2439_adj_1317, n2436_adj_1318, 
        n2435, n2443_adj_1319, n2447_adj_1320, n28228, n2448_adj_1321, 
        n2449_adj_1322, n28319, n2451_adj_1323, n2450_adj_1324, n27964, 
        n2452_adj_1325, n340_adj_1326, n2453_adj_1327, n2454_adj_1328, 
        n38252, n28126, n28420, n1354, n446, n28432, n13606, n14_adj_1332, 
        n4, n26_adj_1333, n2648_adj_1335, n14_adj_1336, n4_adj_1337, 
        n26_adj_1338, n2649_adj_1340, n14_adj_1341, n4_adj_1342, n14_adj_1343, 
        n4_adj_1344, n36747, n20_adj_1345, n6_adj_1346, n2633_adj_1348, 
        n36743, n36760, n36804, n20_adj_1349, n6_adj_1350, n36800, 
        n36817, n36861, n20_adj_1351, n6_adj_1352, n3043_adj_1354, 
        n30740, n2650_adj_1356, n36857, n36874, n3039_adj_1358, n30638, 
        n38293, n591, n2645_adj_1363, n2652_adj_1365, n2642_adj_1367, 
        n2651_adj_1369, n2641_adj_1371, n3052_adj_1373, n36918, n20_adj_1374, 
        n6_adj_1375, n2634_adj_1377, n36914, n36931, n30898, n1845_adj_1379, 
        n3051_adj_1382, n30739, n30738, n30897, n1846_adj_1384, n30637, 
        n3044_adj_1386, n2639_adj_1388, n30636, n30896, n2646_adj_1391, 
        n30895, n38203, n30894, n3047_adj_1398, n2647_adj_1400, n30737, 
        n30893, n30635, n3048_adj_1404, n38208, n12_adj_1406, n28_adj_1407, 
        n30736, n30634, n30735, n30633, n38250, n2654_adj_1413, 
        n2644_adj_1415, n38352, n3032_adj_1417, n2643_adj_1419, n30891, 
        n13638, n28566;
    wire [31:0]n1808_adj_2185;
    
    wire n1743_adj_1421, n1742_adj_1423, n30890, n1745_adj_1425, n38286, 
        n2638_adj_1428, n12429, n38353, n30632, n34948, n30889, 
        n1747_adj_1430, n1746_adj_1432, n2640_adj_1434, n30888, n1749_adj_1436, 
        n1748_adj_1438, n30734, n30631, n30887, n1751_adj_1441, n1750_adj_1443, 
        n30886, n38287, n30732;
    wire [31:0]n2600_adj_2186;
    
    wire n3046_adj_1449, n30629;
    wire [31:0]n1610_adj_2187;
    
    wire n30885, n333_adj_1452, n1754_adj_1454, n30731, n30884, n1643, 
        n30730, n30883, n1645, n38294, n30882, n30881, n38354, 
        n30628, n3035_adj_1469, n30880, n38296, n30879, n3037_adj_1475, 
        n30878, n30729, n30876, n30728, n30875, n38355, n3049_adj_1483, 
        n30727, n30874, n14790, n30873, n30872, n30726, n30725, 
        n36350, n30871, n30724, n30723, n38356, n38357, n30870;
    wire [31:0]n1511;
    
    wire n6_adj_1495, n38408, n38407, n30722, n2537_adj_1498;
    wire [31:0]n2600_adj_2188;
    
    wire n38251, n35636, n28484, n13621;
    wire [31:0]n2897_adj_2189;
    
    wire n2940_adj_1501, n30869, n1745_adj_1502, n35746, n30868, n34788, 
        n5_adj_1503, n38259, n35900, n37596, n37595, n37597, n28267, 
        n13608, n38168, n38213, n12_adj_1506, n28_adj_1507, n3346_adj_1509, 
        n23_adj_1510, n30627, n2951_adj_1514, n30867, n3342_adj_1516, 
        n31_adj_1517, n30626, n3336_adj_1521, n43_adj_1522, n30625, 
        n30866, n30865, n328, n38411, n38181, n3343_adj_1525, n3337_adj_1526, 
        n3332_adj_1527, n38361, n38410, n3128_adj_1528, n34936, n7_adj_1529, 
        n30624, n30721;
    wire [31:0]n2501_adj_2190;
    
    wire n38363, n582, n30623;
    wire [31:0]n1511_adj_2191;
    
    wire n30622, n30863, n30262;
    wire [31:0]n1412_adj_2192;
    
    wire n30720, n10_adj_1540, n38172, n53_adj_1542, n30621, n2932_adj_1546, 
        n349, n3454_adj_1548, n2948_adj_1550, n30240, n38414, n38413, 
        n38365, n2949_adj_1552, n30719, n2934_adj_1556, n3353_adj_1558, 
        n3452_adj_1559, n3334_adj_1561, n47, n13642, n38367, n3351_adj_1563, 
        n13_adj_1564, n10_adj_1565, n2933, n30620, n30619, n3333_adj_1572, 
        n49, n3326_adj_1574, n63_adj_1575, n2936_adj_1577, n2939_adj_1579, 
        n30862, n2930_adj_1583, n38169, n2953_adj_1586, n38170, n2943_adj_1588, 
        n2945_adj_1590, n38417, n2942_adj_1592, n30718, n38266, n38265, 
        n30861, n30860, n38369, n30717, n2442_adj_1601, n30716, 
        n2444_adj_1604, n30715, n38371, n30714, n10_adj_1609, n30859, 
        n30713, n2950_adj_1616, n2938_adj_1618, n2947_adj_1620, n35486, 
        n38416;
    wire [31:0]n2996_adj_2193;
    
    wire n38217, n35142, n38171, n3051_adj_1624, n34720, n28436, 
        n13592, n38210, n38215, n38176, n35302, n35318, n3031_adj_1629, 
        n34904, n30858, n38373, n3045_adj_1633, n30712, n3352, n3353_adj_1636, 
        n3354_adj_1637, n38180, n38058, n38174, n3043_adj_1639, n1742_adj_1640, 
        n3032_adj_1642, n1743_adj_1643, n3040_adj_1645, n30618, n3350_adj_1649, 
        n3046_adj_1651, n3042_adj_1653, n3340_adj_1655, n3035_adj_1657, 
        n38057, n3039_adj_1663, n3030_adj_1665, n3037_adj_1667, n3033_adj_1670, 
        n3036_adj_1673, n3041_adj_1675, n30857, n38298, n3034_adj_1677, 
        n3053_adj_1679, n30856, n30855, n30854, n30852;
    wire [31:0]n1412_adj_2194;
    
    wire n30851, n3054_adj_1686, n30850, n3047_adj_1690, n3048_adj_1692, 
        n3049_adj_1694, n38303, n38301, n3329, n3050_adj_1700, n38218, 
        n30711, n31_adj_1704, n37670, n30709, n13555, n28297;
    wire [31:0]n2402_adj_2195;
    
    wire n2337_adj_1706, n2336_adj_1708, n37504, n3342_adj_1713, n3334_adj_1714, 
        n3345_adj_1715, n3335_adj_1716, n37671, n37515, n36078, n36084, 
        n36074, n36080, n3349_adj_1724, n3129, n3131_adj_1727, n36076, 
        n36056, n3132_adj_1728, n30616, n35780, n28184, n38200, 
        n35462, n35206, n38223, n35466, n348_adj_1735, n3354_adj_1736, 
        n34474, n30708, n2339_adj_1739, n2338_adj_1741, n349_adj_1742, 
        n34078, n30615, n30707, n2341_adj_1744, n2340_adj_1746, n30849, 
        n3340_adj_1749, n34, n37_adj_1750, n339_adj_1752, n596, n34015, 
        n3348_adj_1757, n34013, n35976, n36690, n34594, n588, n38165, 
        n33490, n595, n590, n589, n3232_adj_1767, n38188, n34818, 
        n38375, n30706, n2343, n2342_adj_1771, n10_adj_1772, n30848, 
        n30847;
    wire [31:0]n1511_adj_2196;
    
    wire n3253_adj_1776, n34872, n3230_adj_1779, n30846, n30845, n31270, 
        n13597, n28387, n2139_adj_1785, n2138_adj_1786;
    wire [31:0]n2303_adj_2197;
    
    wire n31269, n2141_adj_1789, n2140_adj_1790, n30614, n31268, n2143_adj_1793, 
        n2142_adj_1794, n31267, n2145_adj_1797, n2144_adj_1798, n30844, 
        n31266, n2147_adj_1803, n2146_adj_1804, n31265, n2149_adj_1807, 
        n2148_adj_1808, n38377, n30705, n2345_adj_1812, n2344_adj_1814, 
        n31264, n2151_adj_1815, n2150_adj_1816, n31263, n2153_adj_1819, 
        n2152_adj_1820, n36698, n36660, n36628, n36630, n36656, 
        n36658, n31262, n2154_adj_1823, n31261, n13616, n28208, 
        n2237_adj_1827;
    wire [31:0]n2402_adj_2198;
    
    wire n30704, n2347_adj_1830, n38270, n31260, n2239_adj_1832, n2238_adj_1833, 
        n31259, n2241_adj_1836, n2240_adj_1837, n31258, n2243_adj_1840, 
        n2242_adj_1841, n31257, n2245_adj_1844, n2244_adj_1845, n31256, 
        n2247_adj_1848, n2246_adj_1849, n31255, n2249_adj_1852, n2248_adj_1853, 
        n31254, n2251_adj_1856, n2250_adj_1857, n30703, n2349_adj_1861, 
        n2348_adj_1863, n30843, n30613, n38381, n38382, n30702, 
        n2351_adj_1867, n2350_adj_1869, n28082, n13601, n30842, n31253, 
        n2253_adj_1872, n2252_adj_1873, n18_adj_1876, n30701, n2353_adj_1878, 
        n2352_adj_1880, n30840;
    wire [31:0]n1610_adj_2199;
    
    wire n30839, n30838, n2540_adj_1888, n31252, n2254_adj_1889, n8_adj_1892, 
        n30837, n30836, n30835, n38383, n30834, n38387, n38388, 
        n31250, n13546, n28022, n38268, n2336_adj_1900;
    wire [31:0]n2501_adj_2200;
    
    wire n18_adj_1903, n30833, n31249, n2339_adj_1904, n2338_adj_1905, 
        n30700, n2354_adj_1910, n30832, n30831, n30830, n30612, 
        n8_adj_1911, n31248, n2341_adj_1912, n2340_adj_1913, n30829, 
        n30699, n13557, n28269, n2237_adj_1916, n30698, n2239_adj_1917, 
        n2238_adj_1918, n38185, n36016, n30828, n38389, n2549_adj_1920, 
        n30697, n2241_adj_1921, n2240_adj_1922, n30826, n30696, n2243_adj_1924, 
        n2242_adj_1925, n38393, n38394, n30825, n2546_adj_1927, n31247, 
        n2343_adj_1928, n2342_adj_1929, n31246, n2345_adj_1932, n2344_adj_1933, 
        n31245, n2347_adj_1936, n2346_adj_1937, n2552_adj_1941, n31244, 
        n2349_adj_1942, n2348_adj_1943, n31243, n2351_adj_1946, n2350_adj_1947, 
        n31242, n2353_adj_1950, n2352_adj_1951, n31241, n2354_adj_1954, 
        n31240, n13599, n28096, n2435_adj_1958, n31239, n38260, 
        n38261, n18_adj_1962, n31238, n2439_adj_1963, n2438_adj_1964, 
        n31237, n2441_adj_1966, n2440, n31236, n2443_adj_1968, n2442_adj_1969, 
        n2534_adj_1972, n31235, n2445_adj_1973, n2444_adj_1974, n31234, 
        n2447_adj_1977, n2446_adj_1978, n31233, n2449_adj_1980, n2448_adj_1981, 
        n31232, n2451_adj_1984, n2450_adj_1985, n31231, n2453_adj_1987, 
        n2452_adj_1988, n31230, n2454_adj_1990, n2539_adj_1993, n31228, 
        n2535_adj_1994, n3147_adj_1996, n34666, n34856, n27858, n8_adj_1997, 
        n2545_adj_1998, n2536_adj_1999, n38256, n38395, n31227, n31226, 
        n2538_adj_2000, n31225, n31224, n2543_adj_2001, n2542_adj_2002, 
        n38399, n38400, n31223, n2544_adj_2003, n31222, n2547_adj_2004, 
        n31221, n2548_adj_2005, n31220, n2551_adj_2006, n2550_adj_2007, 
        n31219, n2553_adj_2008, n31218, n2554_adj_2009, n3148_adj_2011, 
        n18_adj_2012, n8_adj_2013, n31217, n3133_adj_2014, n30695, 
        n2245_adj_2015, n2244_adj_2016, n30824, n36396, n36404, n38253, 
        n36472, n36402, n36470, n36462, n35288, n35294, n35284, 
        n35290, n31216, n31215, n30694, n2247_adj_2017, n2246_adj_2018, 
        n35028, n28303, n13607, n30611, n31214, n31213, n31212, 
        n31211, n28160, n13556, n36654, n31210, n38258, n38257, 
        n35088, n25_adj_2019, n36356, n28_adj_2020, n31209, n31208, 
        n3153_adj_2021, n31207, n31206, n28224, n13619, n35886, 
        n35882, n37672, n37669, n35856, n35854, n35858, n3329_adj_2023, 
        n36022, n3130_adj_2025, n31190, n31189, n31188, n36250, 
        n36246, n36234, n38183, n28237, n27976, n31187, n31186, 
        n31185, n35286, n31184, n3133_adj_2028, n31183, n31182, 
        n31181, n31180, n31179, n31178, n31177, n31176, n31175, 
        n31174, n38206, n31173, n31172, n3138_adj_2031, n31171, 
        n31170, n35790, n35820, n3350_adj_2032, n28172, n3348_adj_2033, 
        n3349_adj_2034, n31169, n31168, n3129_adj_2036, n3140_adj_2038, 
        n38272, n38279, n38284, n38285, n31167, n3145_adj_2040, 
        n36032, n36036, n36026, n36030, n31166, n3128_adj_2042, 
        n34510, n3344_adj_2043, n3328_adj_2044, n3338_adj_2045, n35568, 
        n35566, n3131_adj_2047, n38167, n3333_adj_2048, n31164, n31163, 
        n31162, n31161, n28158, n31160, n31159, n31158, n27882, 
        n31157, n31156, n3144_adj_2067, n38264, n35590, n31155, 
        n35588, n38263, n3134_adj_2070, n35584, n35582, n31154, 
        n28154, n27876, n3146_adj_2073, n35902, n35898, n3141_adj_2075, 
        n30823, n31153, n31152, n30822, n35940, n38418, n35938, 
        n3139_adj_2080, n30821, n38267, n30610, n34956, n34958, 
        n31151, n31150, n31149, n31148, n31147, n35534, n35526, 
        n35532, n31146, n31145, n31144, n27996, n27745, n36264, 
        n36262, n31143, n31142, n28241, n2248_adj_2086, n2249_adj_2087, 
        n31141, n2251_adj_2089, n2250_adj_2090, n27982, n2252_adj_2091, 
        n2253_adj_2092, n2254_adj_2093, n35606, n31140, n35602, n27988, 
        n27735, n35096, n35060, n3137_adj_2096, n35092, n3136_adj_2097, 
        n27970, n31139, n31138, n27199, n3142_adj_2101, n38204, 
        n35648, n35642, n35644, n34804, n5_adj_2103, n27994, n27749, 
        n28192, n27923, n37517, n35130, n35132, n37506, n35102, 
        n35106, n37488, n35110, n3154_adj_2106, n31136, n31135, 
        n35498, n35496, n33697, n35494, n28289, n28040, n31134, 
        n35394, n35392, n35390, n31133, n31132, n31131, n28279, 
        n28506, n28024, n2952_adj_2110, n345_adj_2111, n2954_adj_2112, 
        n35262, n35252, n13618, n35260, n31130, n31129, n2937_adj_2113, 
        n2935_adj_2114, n35254, n35240, n34912, n28002, n30820, 
        n35334, n35330, n35322, n35324, n35328, n2931_adj_2115, 
        n2946_adj_2116, n2944_adj_2117, n31128, n31127, n28285, n28030, 
        n344_adj_2118, n31126, n3149_adj_2119, n31125, n3150_adj_2120, 
        n35468, n35476, n35472, n38205, n28271, n28014, n35368, 
        n35366, n35362, n35358, n28277, n28018, n35050, n35000, 
        n34998, n34988, n35046, n35042, n31124, n31123, n37668, 
        n28261, n28010, n31122, n35036, n35020, n35016, n35018, 
        n35032, n31121, n31120, n31119, n36650, n36899, n36886, 
        n5_adj_2121, n31118, n31117, n36842, n33434, n36829, n31116, 
        n34880, n34790, n28098, n5_adj_2122, n31115, n36785, n35728, 
        n36772, n5_adj_2123, n36728, n36715, n5_adj_2124, n31114, 
        n31113, n28391, n28110, n31112, n38269;
    wire [31:0]n2996_adj_2201;
    
    wire n38209, n31539, n34944, n34942, n31111, n31110, n31109, 
        n31108, n31107, n31106, n31105, n31104, n31103, n31101, 
        n31100, n31099, n38271, n36316, n36318, n36310, n36314, 
        n35930, n35784, n27984, n31098, n31097, n38166, n31096, 
        n31095, n31094, n31093, n31092, n31091, n31090, n31089, 
        n31088, n31087, n31086, n31085, n31084, n31083, n31082, 
        n31081, n34774, n34772, n31080, n31079, n31078, n31077, 
        n31075, n31074, n31073, n31072, n31071, n31070, n31069, 
        n31068, n31067, n31066, n31065, n31064, n31063, n31062, 
        n31061, n31060, n31059, n31058, n31057, n31056, n31055, 
        n31054, n31052, n31051, n31050, n31049, n31048, n31047, 
        n31046, n31045, n31044, n31043, n38276, n31042, n31041, 
        n31040, n31039, n38207, n34812, n31038, n31037, n35176, 
        n31036, n31035, n35082, n35068, n35078, n28293, n28042, 
        n31034, n31033, n31032, n31031, n31030, n31029, n31028, 
        n31027, n31026, n34766, n27919, n31025, n31023, n34836, 
        n33591, n31022, n31021, n34852, n34710, n34928, n27862, 
        n35192, n35198, n35188, n35194, n35190, n34700, n27878, 
        n35162, n35164, n35156, n35160, n31020, n31019, n31018, 
        n35150, n31017, n31016, n31015, n31014, n31013, n31012, 
        n34810, n27888, n35226, n35228, n35220, n35224, n31011, 
        n34658, n27905, n35440, n35448, n35444, n31010, n31009, 
        n34728, n27915, n35420, n35418, n35416, n31008, n31007, 
        n31006, n31005, n31004, n31003, n31002, n31001, n31000, 
        n30999, n30998, n38288, n38214, n34129, n34970, n30996, 
        n30995, n34966, n10_adj_2159, n30819, n30818, n30817, n30994, 
        n30693, n30993, n30692, n30816, n30815, n30992, n30991, 
        n30691, n30813, n30990, n30989, n30988, n30690, n30987, 
        n30986, n30985, n30984, n30983, n30812, n30982, n30981;
    
    LUT4 i1_2_lut_4_lut (.A(n1744), .B(n1808[29]), .C(n38295), .D(n1846), 
         .Z(n35744)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut.init = 16'hffca;
    CCU2C rem_10_add_1244_11 (.A0(n13631), .B0(n28090), .C0(n1808[25]), 
          .D0(n1748), .A1(n13631), .B1(n28090), .C1(n1808[26]), .D1(n1747), 
          .CIN(n30608), .COUT(n30609), .S0(n1907[25]), .S1(n1907[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_11.INIT0 = 16'hf1e0;
    defparam rem_10_add_1244_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1244_11.INJECT1_0 = "NO";
    defparam rem_10_add_1244_11.INJECT1_1 = "NO";
    CCU2C div_9_add_2182_23 (.A0(n13547), .B0(n28588), .C0(n3194[24]), 
          .D0(n3135), .A1(n13547), .B1(n28588), .C1(n3194[25]), .D1(n3134), 
          .CIN(n30810), .COUT(n30811), .S0(n3293[24]), .S1(n3293[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_23.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_23.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_23.INJECT1_0 = "NO";
    defparam div_9_add_2182_23.INJECT1_1 = "NO";
    LUT4 i26566_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[27]), 
         .D(n2[19]), .Z(n1746)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26566_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1917_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[30]), 
         .D(n2832), .Z(n2931)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1917_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i26531_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[29]), 
         .D(n35[19]), .Z(n1744_adj_520)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26531_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1933_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[14]), 
         .D(n2848), .Z(n2947)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1933_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1244_9 (.A0(n13631), .B0(n28090), .C0(n1808[23]), 
          .D0(n1750), .A1(n13631), .B1(n28090), .C1(n1808[24]), .D1(n1749), 
          .CIN(n30607), .COUT(n30608), .S0(n1907[23]), .S1(n1907[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1244_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1244_9.INJECT1_0 = "NO";
    defparam rem_10_add_1244_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1244_7 (.A0(n13631), .B0(n28090), .C0(n1808[21]), 
          .D0(n1752), .A1(n13631), .B1(n28090), .C1(n1808[22]), .D1(n1751), 
          .CIN(n30606), .COUT(n30607), .S0(n1907[21]), .S1(n1907[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_7.INIT0 = 16'hf1e0;
    defparam rem_10_add_1244_7.INIT1 = 16'h0e1f;
    defparam rem_10_add_1244_7.INJECT1_0 = "NO";
    defparam rem_10_add_1244_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1512_19 (.A0(n13590), .B0(n28440), .C0(n2204[30]), 
          .D0(n38275), .A1(n13590), .B1(n28440), .C1(n2204[31]), .D1(n38274), 
          .CIN(n30688), .S0(n2303[30]), .S1(n2303[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1512_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1512_19.INJECT1_0 = "NO";
    defparam div_9_add_1512_19.INJECT1_1 = "NO";
    FD1S3IX pwm_cnt_1138__i0 (.D(n50[0]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i0.GSR = "ENABLED";
    LUT4 div_9_i1923_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[24]), 
         .D(n2838), .Z(n2937)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1923_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2198_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[17]), 
         .D(n3241), .Z(n3340)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2198_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_26227_31 (.A0(n13629), .B0(n28492), .C0(n3293[31]), .D0(n3227), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n30547), 
          .S0(n3392[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_31.INIT0 = 16'h0e1f;
    defparam add_26227_31.INIT1 = 16'h0000;
    defparam add_26227_31.INJECT1_0 = "NO";
    defparam add_26227_31.INJECT1_1 = "NO";
    LUT4 rem_10_i2203_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[12]), 
         .D(n3246), .Z(n3345)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2203_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_26227_29 (.A0(n13629), .B0(n28492), .C0(n3293[29]), .D0(n38190), 
          .A1(n13629), .B1(n28492), .C1(n3293[30]), .D1(n3228), .CIN(n30546), 
          .COUT(n30547), .S0(n3392[29]), .S1(n3392[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_29.INIT0 = 16'h0e1f;
    defparam add_26227_29.INIT1 = 16'h0e1f;
    defparam add_26227_29.INJECT1_0 = "NO";
    defparam add_26227_29.INJECT1_1 = "NO";
    CCU2C rem_10_add_1244_5 (.A0(n13631), .B0(n28090), .C0(n1808[19]), 
          .D0(n1754), .A1(n13631), .B1(n28090), .C1(n1808[20]), .D1(n1753), 
          .CIN(n30605), .COUT(n30606), .S0(n1907[19]), .S1(n1907[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_5.INIT0 = 16'h0e1f;
    defparam rem_10_add_1244_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1244_5.INJECT1_0 = "NO";
    defparam rem_10_add_1244_5.INJECT1_1 = "NO";
    LUT4 rem_10_i2367_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[6]), .D(n3549), 
         .Z(n36[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2367_3_lut_4_lut.init = 16'hf780;
    CCU2C rem_10_add_1244_3 (.A0(n12154), .B0(n5), .C0(n39), .D0(n2[17]), 
          .A1(n38307), .B1(n1808[18]), .C1(n2[18]), .D1(n38295), .CIN(n30604), 
          .COUT(n30605), .S0(n1907[17]), .S1(n1907[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_3.INIT0 = 16'h5410;
    defparam rem_10_add_1244_3.INIT1 = 16'hcca0;
    defparam rem_10_add_1244_3.INJECT1_0 = "NO";
    defparam rem_10_add_1244_3.INJECT1_1 = "NO";
    CCU2C div_9_add_1512_17 (.A0(n13590), .B0(n28440), .C0(n2204[28]), 
          .D0(n2141), .A1(n13590), .B1(n28440), .C1(n2204[29]), .D1(n2140), 
          .CIN(n30687), .COUT(n30688), .S0(n2303[28]), .S1(n2303[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1512_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1512_17.INJECT1_0 = "NO";
    defparam div_9_add_1512_17.INJECT1_1 = "NO";
    LUT4 rem_10_mux_3_i7_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[6]), .D(duty0_14__N_426[4]), 
         .Z(n594)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i7_3_lut_4_lut.init = 16'hf780;
    CCU2C div_9_add_2182_21 (.A0(n13547), .B0(n28588), .C0(n3194[22]), 
          .D0(n3137), .A1(n13547), .B1(n28588), .C1(n3194[23]), .D1(n3136), 
          .CIN(n30809), .COUT(n30810), .S0(n3293[22]), .S1(n3293[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_21.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_21.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_21.INJECT1_0 = "NO";
    defparam div_9_add_2182_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_11 (.A(n2853), .B(n2897_adj_2162[9]), .C(n38226), 
         .D(n2951), .Z(n34692)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_11.init = 16'hca00;
    LUT4 rem_10_i2190_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[25]), 
         .D(n3233), .Z(n3332)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2190_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2182_19 (.A0(n13547), .B0(n28588), .C0(n3194[20]), 
          .D0(n3139), .A1(n13547), .B1(n28588), .C1(n3194[21]), .D1(n3138), 
          .CIN(n30808), .COUT(n30809), .S0(n3293[20]), .S1(n3293[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_19.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_19.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_19.INJECT1_0 = "NO";
    defparam div_9_add_2182_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_12 (.A(n2842), .B(n2897_adj_2162[20]), .C(n38226), 
         .D(n2940), .Z(n35208)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_12.init = 16'hffca;
    LUT4 rem_10_i2365_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[8]), .D(n3547), 
         .Z(n36[8])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2365_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i2366_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[7]), .D(n3548), 
         .Z(n36[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2366_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_mux_3_i14_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[13]), 
         .D(duty0_14__N_426[11]), .Z(n587)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 i24430_2_lut_rep_221 (.A(n28307), .B(n13598), .Z(n38226)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24430_2_lut_rep_221.init = 16'heeee;
    LUT4 i1_3_lut (.A(n27382), .B(n3), .C(distance[0]), .Z(duty0_14__N_426[0])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h2020;
    LUT4 rem_10_i1919_3_lut_rep_215_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[28]), 
         .D(n2834), .Z(n38220)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1919_3_lut_rep_215_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1938_3_lut_rep_219_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[9]), 
         .D(n2853), .Z(n38224)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1938_3_lut_rep_219_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2368_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[5]), .D(n3550), 
         .Z(n36[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2368_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i1927_3_lut_rep_220_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[20]), 
         .D(n2842), .Z(n38225)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1927_3_lut_rep_220_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2364_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[9]), .D(n3546), 
         .Z(n36[9])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2364_3_lut_4_lut.init = 16'hf780;
    CCU2C add_26227_27 (.A0(n13629), .B0(n28492), .C0(n3293[27]), .D0(n3231), 
          .A1(n13629), .B1(n28492), .C1(n3293[28]), .D1(n3230), .CIN(n30545), 
          .COUT(n30546), .S0(n3392[27]), .S1(n3392[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_27.INIT0 = 16'h0e1f;
    defparam add_26227_27.INIT1 = 16'h0e1f;
    defparam add_26227_27.INJECT1_0 = "NO";
    defparam add_26227_27.INJECT1_1 = "NO";
    FD1S3JX duty0_i0 (.D(duty0_14__N_410[0]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i0.GSR = "DISABLED";
    LUT4 rem_10_i2371_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[2]), .D(n3454), 
         .Z(n36[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2371_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i2369_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[4]), .D(n3551), 
         .Z(n36[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2369_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i2341_4_lut (.A(n38179), .B(n3449), .C(n3458), .D(n38175), 
         .Z(n3547)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2341_4_lut.init = 16'h6aaa;
    CCU2C add_26227_25 (.A0(n13629), .B0(n28492), .C0(n3293[25]), .D0(n3233_adj_522), 
          .A1(n13629), .B1(n28492), .C1(n3293[26]), .D1(n3232), .CIN(n30544), 
          .COUT(n30545), .S0(n3392[25]), .S1(n3392[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_25.INIT0 = 16'h0e1f;
    defparam add_26227_25.INIT1 = 16'h0e1f;
    defparam add_26227_25.INJECT1_0 = "NO";
    defparam add_26227_25.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n34756), .B(n33580), .C(n34758), .D(n39_adj_523), 
         .Z(n3458)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 rem_10_i1916_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[31]), 
         .D(n38229), .Z(n2930)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1916_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1244_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n42), .D1(n2[16]), 
          .COUT(n30604));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_1.INIT0 = 16'h000F;
    defparam rem_10_add_1244_1.INIT1 = 16'habef;
    defparam rem_10_add_1244_1.INJECT1_0 = "NO";
    defparam rem_10_add_1244_1.INJECT1_1 = "NO";
    FD1S3JX duty1_i0 (.D(duty1_14__N_458[0]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i0.GSR = "DISABLED";
    FD1S3JX duty2_i0 (.D(duty2_14__N_473[0]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i0.GSR = "DISABLED";
    FD1S3JX duty3_i0 (.D(duty3_14__N_488[0]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i0.GSR = "DISABLED";
    CCU2C div_9_add_909_11 (.A0(n27382), .B0(n3), .C0(n5), .D0(n35[19]), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n30603), 
          .S0(n1412[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_909_11.INIT0 = 16'hffff;
    defparam div_9_add_909_11.INIT1 = 16'h0000;
    defparam div_9_add_909_11.INJECT1_0 = "NO";
    defparam div_9_add_909_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1512_15 (.A0(n13590), .B0(n28440), .C0(n2204[26]), 
          .D0(n2143), .A1(n13590), .B1(n28440), .C1(n2204[27]), .D1(n2142), 
          .CIN(n30686), .COUT(n30687), .S0(n2303[26]), .S1(n2303[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1512_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1512_15.INJECT1_0 = "NO";
    defparam div_9_add_1512_15.INJECT1_1 = "NO";
    CCU2C add_26227_23 (.A0(n13629), .B0(n28492), .C0(n3293[23]), .D0(n3235), 
          .A1(n13629), .B1(n28492), .C1(n3293[24]), .D1(n3234), .CIN(n30543), 
          .COUT(n30544), .S0(n3392[23]), .S1(n3392[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_23.INIT0 = 16'h0e1f;
    defparam add_26227_23.INIT1 = 16'h0e1f;
    defparam add_26227_23.INJECT1_0 = "NO";
    defparam add_26227_23.INJECT1_1 = "NO";
    CCU2C div_9_add_909_9 (.A0(n27382), .B0(n3), .C0(n5), .D0(n35[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), .CIN(n30602), 
          .COUT(n30603), .S0(n1412[29]), .S1(n1412[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_909_9.INIT0 = 16'h0000;
    defparam div_9_add_909_9.INIT1 = 16'h0000;
    defparam div_9_add_909_9.INJECT1_0 = "NO";
    defparam div_9_add_909_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_13 (.A(n3435), .B(n34752), .C(n34740), .D(n3437), 
         .Z(n34756)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_13.init = 16'hfffe;
    LUT4 rem_10_i1923_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[24]), 
         .D(n2838_adj_525), .Z(n2937_adj_526)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1923_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_mux_3_i15_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[14]), 
         .D(duty0_14__N_426[12]), .Z(n586)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i1928_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[19]), 
         .D(n2843), .Z(n2942)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1928_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_14 (.A(n3446), .B(n31), .C(n34746), .D(n3434), 
         .Z(n34758)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_14.init = 16'hfffe;
    CCU2C div_9_add_2182_17 (.A0(n13547), .B0(n28588), .C0(n3194[18]), 
          .D0(n3141), .A1(n13547), .B1(n28588), .C1(n3194[19]), .D1(n3140), 
          .CIN(n30807), .COUT(n30808), .S0(n3293[18]), .S1(n3293[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_17.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_17.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_17.INJECT1_0 = "NO";
    defparam div_9_add_2182_17.INJECT1_1 = "NO";
    CCU2C div_9_add_2182_15 (.A0(n13547), .B0(n28588), .C0(n3194[16]), 
          .D0(n38201), .A1(n13547), .B1(n28588), .C1(n3194[17]), .D1(n3142), 
          .CIN(n30806), .COUT(n30807), .S0(n3293[16]), .S1(n3293[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_15.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_15.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_15.INJECT1_0 = "NO";
    defparam div_9_add_2182_15.INJECT1_1 = "NO";
    CCU2C div_13_add_1847_15 (.A0(n13624), .B0(n28462), .C0(n2699[21]), 
          .D0(n2643), .A1(n13624), .B1(n28462), .C1(n2699[22]), .D1(n2642), 
          .CIN(n30979), .COUT(n30980), .S0(n2798[21]), .S1(n2798[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_15.INJECT1_0 = "NO";
    defparam div_13_add_1847_15.INJECT1_1 = "NO";
    LUT4 i26572_3_lut_4_lut (.A(n5), .B(n38331), .C(n4540[20]), .D(n4540[18]), 
         .Z(n31386)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26572_3_lut_4_lut.init = 16'h8880;
    LUT4 i1_4_lut_adj_15 (.A(n3443), .B(n3440), .C(n3436), .D(n3441), 
         .Z(n34752)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_15.init = 16'hfffe;
    LUT4 mux_1857_i6_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[7]), .D(duty0_14__N_426[5]), 
         .Z(n344)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i6_3_lut_4_lut.init = 16'hf780;
    CCU2C div_13_add_1847_13 (.A0(n13624), .B0(n28462), .C0(n2699[19]), 
          .D0(n2645), .A1(n13624), .B1(n28462), .C1(n2699[20]), .D1(n2644), 
          .CIN(n30978), .COUT(n30979), .S0(n2798[19]), .S1(n2798[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_13.INJECT1_0 = "NO";
    defparam div_13_add_1847_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1925_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[22]), 
         .D(n38238), .Z(n2939)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1925_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1857_i16_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[17]), .D(duty0_14__N_426[15]), 
         .Z(n334)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i1932_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[15]), 
         .D(n2847), .Z(n2946)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1932_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1857_i12_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[13]), .D(duty0_14__N_426[11]), 
         .Z(n338)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i12_3_lut_4_lut.init = 16'hf780;
    CCU2C div_13_add_1847_11 (.A0(n13624), .B0(n28462), .C0(n2699[17]), 
          .D0(n2647), .A1(n13624), .B1(n28462), .C1(n2699[18]), .D1(n2646), 
          .CIN(n30977), .COUT(n30978), .S0(n2798[17]), .S1(n2798[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_11.INJECT1_0 = "NO";
    defparam div_13_add_1847_11.INJECT1_1 = "NO";
    LUT4 rem_10_i2276_3_lut (.A(n3351), .B(n3392_adj_2163[6]), .C(n3359), 
         .Z(n3450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2276_3_lut.init = 16'hcaca;
    CCU2C div_13_add_1847_9 (.A0(n13624), .B0(n28462), .C0(n2699[15]), 
          .D0(n2649), .A1(n13624), .B1(n28462), .C1(n2699[16]), .D1(n2648), 
          .CIN(n30976), .COUT(n30977), .S0(n2798[15]), .S1(n2798[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1847_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1847_9.INJECT1_0 = "NO";
    defparam div_13_add_1847_9.INJECT1_1 = "NO";
    CCU2C div_9_add_909_7 (.A0(n27382), .B0(n3), .C0(n5), .D0(n35[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), .CIN(n30601), 
          .COUT(n30602), .S0(n1412[27]), .S1(n1412[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_909_7.INIT0 = 16'hffff;
    defparam div_9_add_909_7.INIT1 = 16'h2000;
    defparam div_9_add_909_7.INJECT1_0 = "NO";
    defparam div_9_add_909_7.INJECT1_1 = "NO";
    LUT4 mux_1857_i5_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[6]), .D(duty0_14__N_426[4]), 
         .Z(n345)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i5_3_lut_4_lut.init = 16'hf780;
    CCU2C div_9_add_1512_13 (.A0(n13590), .B0(n28440), .C0(n2204[24]), 
          .D0(n38277), .A1(n13590), .B1(n28440), .C1(n2204[25]), .D1(n2144), 
          .CIN(n30685), .COUT(n30686), .S0(n2303[24]), .S1(n2303[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1512_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1512_13.INJECT1_0 = "NO";
    defparam div_9_add_1512_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1924_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[23]), 
         .D(n2839), .Z(n2938)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1924_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2182_13 (.A0(n13547), .B0(n28588), .C0(n3194[14]), 
          .D0(n3145), .A1(n13547), .B1(n28588), .C1(n3194[15]), .D1(n3144), 
          .CIN(n30805), .COUT(n30806), .S0(n3293[14]), .S1(n3293[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_13.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_13.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_13.INJECT1_0 = "NO";
    defparam div_9_add_2182_13.INJECT1_1 = "NO";
    CCU2C div_9_add_2182_11 (.A0(n13547), .B0(n28588), .C0(n3194[12]), 
          .D0(n3147), .A1(n13547), .B1(n28588), .C1(n3194[13]), .D1(n3146), 
          .CIN(n30804), .COUT(n30805), .S0(n3293[12]), .S1(n3293[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_11.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_11.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_11.INJECT1_0 = "NO";
    defparam div_9_add_2182_11.INJECT1_1 = "NO";
    CCU2C div_13_add_1847_7 (.A0(n13624), .B0(n28462), .C0(n2699[13]), 
          .D0(n2651), .A1(n13624), .B1(n28462), .C1(n2699[14]), .D1(n2650), 
          .CIN(n30975), .COUT(n30976), .S0(n2798[13]), .S1(n2798[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1847_7.INJECT1_0 = "NO";
    defparam div_13_add_1847_7.INJECT1_1 = "NO";
    LUT4 rem_10_mux_3_i16_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[15]), 
         .D(duty0_14__N_426[13]), .Z(n585)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1857_i9_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[10]), .D(duty0_14__N_426[8]), 
         .Z(n341)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_i2278_3_lut (.A(n3353), .B(n3392_adj_2163[4]), .C(n3359), 
         .Z(n3452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2278_3_lut.init = 16'hcaca;
    CCU2C div_9_add_1512_11 (.A0(n13590), .B0(n28440), .C0(n2204[22]), 
          .D0(n2147), .A1(n13590), .B1(n28440), .C1(n2204[23]), .D1(n2146), 
          .CIN(n30684), .COUT(n30685), .S0(n2303[22]), .S1(n2303[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1512_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1512_11.INJECT1_0 = "NO";
    defparam div_9_add_1512_11.INJECT1_1 = "NO";
    CCU2C add_26227_21 (.A0(n13629), .B0(n28492), .C0(n3293[21]), .D0(n3237), 
          .A1(n13629), .B1(n28492), .C1(n3293[22]), .D1(n3236), .CIN(n30542), 
          .COUT(n30543), .S0(n3392[21]), .S1(n3392[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_21.INIT0 = 16'h0e1f;
    defparam add_26227_21.INIT1 = 16'h0e1f;
    defparam add_26227_21.INJECT1_0 = "NO";
    defparam add_26227_21.INJECT1_1 = "NO";
    CCU2C add_26227_19 (.A0(n13629), .B0(n28492), .C0(n3293[19]), .D0(n3239), 
          .A1(n13629), .B1(n28492), .C1(n3293[20]), .D1(n3238), .CIN(n30541), 
          .COUT(n30542), .S0(n3392[19]), .S1(n3392[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_19.INIT0 = 16'h0e1f;
    defparam add_26227_19.INIT1 = 16'h0e1f;
    defparam add_26227_19.INJECT1_0 = "NO";
    defparam add_26227_19.INJECT1_1 = "NO";
    LUT4 rem_10_i1926_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[21]), 
         .D(n2841), .Z(n2940)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1926_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_909_5 (.A0(n27382), .B0(n3), .C0(n5), .D0(n35[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), .CIN(n30600), 
          .COUT(n30601), .S0(n1412[25]), .S1(n1412[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_909_5.INIT0 = 16'h2000;
    defparam div_9_add_909_5.INIT1 = 16'h0000;
    defparam div_9_add_909_5.INJECT1_0 = "NO";
    defparam div_9_add_909_5.INJECT1_1 = "NO";
    CCU2C add_26227_17 (.A0(n13629), .B0(n28492), .C0(n3293[17]), .D0(n3241_adj_532), 
          .A1(n13629), .B1(n28492), .C1(n3293[18]), .D1(n3240), .CIN(n30540), 
          .COUT(n30541), .S0(n3392[17]), .S1(n3392[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_17.INIT0 = 16'h0e1f;
    defparam add_26227_17.INIT1 = 16'h0e1f;
    defparam add_26227_17.INJECT1_0 = "NO";
    defparam add_26227_17.INJECT1_1 = "NO";
    CCU2C add_26227_15 (.A0(n13629), .B0(n28492), .C0(n3293[15]), .D0(n3243), 
          .A1(n13629), .B1(n28492), .C1(n3293[16]), .D1(n3242), .CIN(n30539), 
          .COUT(n30540), .S0(n3392[15]), .S1(n3392[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_15.INIT0 = 16'h0e1f;
    defparam add_26227_15.INIT1 = 16'h0e1f;
    defparam add_26227_15.INJECT1_0 = "NO";
    defparam add_26227_15.INJECT1_1 = "NO";
    LUT4 rem_10_i1939_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[8]), 
         .D(n2854), .Z(n2953)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1939_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2279_3_lut (.A(n3354), .B(n3392_adj_2163[3]), .C(n3359), 
         .Z(n3453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2279_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1920_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[27]), 
         .D(n2835), .Z(n2934)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1920_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1917_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[30]), 
         .D(n2832_adj_534), .Z(n2931_adj_535)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1917_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_909_3 (.A0(n27382), .B0(n3), .C0(n5), .D0(n35[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), .CIN(n30599), 
          .COUT(n30600), .S0(n1412[23]), .S1(n1412[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_909_3.INIT0 = 16'h0000;
    defparam div_9_add_909_3.INIT1 = 16'hffff;
    defparam div_9_add_909_3.INJECT1_0 = "NO";
    defparam div_9_add_909_3.INJECT1_1 = "NO";
    CCU2C div_9_add_909_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), .COUT(n30599), 
          .S1(n1412[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_909_1.INIT0 = 16'h0000;
    defparam div_9_add_909_1.INIT1 = 16'hdfff;
    defparam div_9_add_909_1.INJECT1_0 = "NO";
    defparam div_9_add_909_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1512_9 (.A0(n13590), .B0(n28440), .C0(n2204[20]), 
          .D0(n2149), .A1(n13590), .B1(n28440), .C1(n2204[21]), .D1(n2148), 
          .CIN(n30683), .COUT(n30684), .S0(n2303[20]), .S1(n2303[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1512_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1512_9.INJECT1_0 = "NO";
    defparam div_9_add_1512_9.INJECT1_1 = "NO";
    LUT4 rem_10_i2277_3_lut (.A(n38187), .B(n3392_adj_2163[5]), .C(n3359), 
         .Z(n3451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2277_3_lut.init = 16'hcaca;
    PFUMX i32314 (.BLUT(n37665), .ALUT(n37664), .C0(n38177), .Z(n37666));
    CCU2C rem_10_add_1311_17 (.A0(n13600), .B0(n28359), .C0(n1907[30]), 
          .D0(n1842), .A1(n13600), .B1(n28359), .C1(n1907[31]), .D1(n1841), 
          .CIN(n30597), .S0(n2006[30]), .S1(n2006[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1311_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1311_17.INJECT1_0 = "NO";
    defparam rem_10_add_1311_17.INJECT1_1 = "NO";
    LUT4 rem_10_i2259_3_lut (.A(n3334), .B(n3392_adj_2163[23]), .C(n3359), 
         .Z(n3433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2259_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2207_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[8]), 
         .D(n3250), .Z(n3349)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2207_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2188_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[27]), 
         .D(n38191), .Z(n3330)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1921_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[26]), 
         .D(n2836), .Z(n2935)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1921_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2192_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[23]), 
         .D(n3235_adj_539), .Z(n3334)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2192_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_26227_13 (.A0(n13629), .B0(n28492), .C0(n3293[13]), .D0(n3245), 
          .A1(n13629), .B1(n28492), .C1(n3293[14]), .D1(n3244), .CIN(n30538), 
          .COUT(n30539), .S0(n3392[13]), .S1(n3392[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_13.INIT0 = 16'h0e1f;
    defparam add_26227_13.INIT1 = 16'h0e1f;
    defparam add_26227_13.INJECT1_0 = "NO";
    defparam add_26227_13.INJECT1_1 = "NO";
    LUT4 rem_10_i2272_3_lut (.A(n3347), .B(n3392_adj_2163[10]), .C(n3359), 
         .Z(n3446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2272_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1930_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[17]), 
         .D(n2845), .Z(n2944)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1930_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10_4_lut (.A(n3346), .B(n3438), .C(n3392_adj_2163[11]), .D(n3359), 
         .Z(n31)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i10_4_lut.init = 16'hfcee;
    LUT4 rem_10_i2264_3_lut (.A(n3339), .B(n3392_adj_2163[18]), .C(n3359), 
         .Z(n3438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2264_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1929_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[18]), 
         .D(n2844), .Z(n2943)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1929_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2194_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[21]), 
         .D(n3237_adj_542), .Z(n3336)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2194_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2260_3_lut (.A(n3335), .B(n3392_adj_2163[22]), .C(n3359), 
         .Z(n3434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2260_3_lut.init = 16'hcaca;
    MULT18X18D mult_11_mult_2 (.A17(n36[10]), .A16(n36[10]), .A15(n36[10]), 
            .A14(n36[10]), .A13(n36[10]), .A12(n36[10]), .A11(n36[10]), 
            .A10(n36[10]), .A9(n36[9]), .A8(n36[8]), .A7(n36[7]), .A6(n36[6]), 
            .A5(n36[5]), .A4(n36[4]), .A3(n36[3]), .A2(n36[2]), .A1(n36[1]), 
            .A0(GND_net), .B17(GND_net), .B16(GND_net), .B15(GND_net), 
            .B14(VCC_net), .B13(VCC_net), .B12(GND_net), .B11(GND_net), 
            .B10(GND_net), .B9(GND_net), .B8(VCC_net), .B7(VCC_net), 
            .B6(GND_net), .B5(VCC_net), .B4(GND_net), .B3(GND_net), 
            .B2(VCC_net), .B1(VCC_net), .B0(VCC_net), .C17(GND_net), 
            .C16(GND_net), .C15(GND_net), .C14(GND_net), .C13(GND_net), 
            .C12(GND_net), .C11(GND_net), .C10(GND_net), .C9(GND_net), 
            .C8(GND_net), .C7(GND_net), .C6(GND_net), .C5(GND_net), 
            .C4(GND_net), .C3(GND_net), .C2(GND_net), .C1(GND_net), 
            .C0(GND_net), .SIGNEDA(VCC_net), .SIGNEDB(VCC_net), .SOURCEA(GND_net), 
            .SOURCEB(GND_net), .CLK3(GND_net), .CLK2(GND_net), .CLK1(GND_net), 
            .CLK0(GND_net), .CE3(GND_net), .CE2(GND_net), .CE1(GND_net), 
            .CE0(VCC_net), .RST3(GND_net), .RST2(GND_net), .RST1(GND_net), 
            .RST0(GND_net), .SRIA17(GND_net), .SRIA16(GND_net), .SRIA15(GND_net), 
            .SRIA14(GND_net), .SRIA13(GND_net), .SRIA12(GND_net), .SRIA11(GND_net), 
            .SRIA10(GND_net), .SRIA9(GND_net), .SRIA8(GND_net), .SRIA7(GND_net), 
            .SRIA6(GND_net), .SRIA5(GND_net), .SRIA4(GND_net), .SRIA3(GND_net), 
            .SRIA2(GND_net), .SRIA1(GND_net), .SRIA0(GND_net), .SRIB17(GND_net), 
            .SRIB16(GND_net), .SRIB15(GND_net), .SRIB14(GND_net), .SRIB13(GND_net), 
            .SRIB12(GND_net), .SRIB11(GND_net), .SRIB10(GND_net), .SRIB9(GND_net), 
            .SRIB8(GND_net), .SRIB7(GND_net), .SRIB6(GND_net), .SRIB5(GND_net), 
            .SRIB4(GND_net), .SRIB3(GND_net), .SRIB2(GND_net), .SRIB1(GND_net), 
            .SRIB0(GND_net), .P26(n136), .P25(n58), .P24(n59), .P23(n60), 
            .P22(n61), .P21(n62), .P20(n63), .P19(n64), .P18(n65), 
            .P17(n66), .P16(n67), .P15(n68), .P14(n69), .P13(n70), 
            .P12(n71), .P11(n72), .P10(n73), .P9(n74), .P8(n75), .P7(n76), 
            .P6(n77), .P5(n78), .P4(n79), .P3(n80), .P2(n81), .P1(n82), 
            .P0(n83));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(74[17:32])
    defparam mult_11_mult_2.REG_INPUTA_CLK = "NONE";
    defparam mult_11_mult_2.REG_INPUTA_CE = "CE0";
    defparam mult_11_mult_2.REG_INPUTA_RST = "RST0";
    defparam mult_11_mult_2.REG_INPUTB_CLK = "NONE";
    defparam mult_11_mult_2.REG_INPUTB_CE = "CE0";
    defparam mult_11_mult_2.REG_INPUTB_RST = "RST0";
    defparam mult_11_mult_2.REG_INPUTC_CLK = "NONE";
    defparam mult_11_mult_2.REG_INPUTC_CE = "CE0";
    defparam mult_11_mult_2.REG_INPUTC_RST = "RST0";
    defparam mult_11_mult_2.REG_PIPELINE_CLK = "NONE";
    defparam mult_11_mult_2.REG_PIPELINE_CE = "CE0";
    defparam mult_11_mult_2.REG_PIPELINE_RST = "RST0";
    defparam mult_11_mult_2.REG_OUTPUT_CLK = "NONE";
    defparam mult_11_mult_2.REG_OUTPUT_CE = "CE0";
    defparam mult_11_mult_2.REG_OUTPUT_RST = "RST0";
    defparam mult_11_mult_2.CLK0_DIV = "ENABLED";
    defparam mult_11_mult_2.CLK1_DIV = "ENABLED";
    defparam mult_11_mult_2.CLK2_DIV = "ENABLED";
    defparam mult_11_mult_2.CLK3_DIV = "ENABLED";
    defparam mult_11_mult_2.HIGHSPEED_CLK = "NONE";
    defparam mult_11_mult_2.GSR = "DISABLED";
    defparam mult_11_mult_2.CAS_MATCH_REG = "FALSE";
    defparam mult_11_mult_2.SOURCEB_MODE = "B_SHIFT";
    defparam mult_11_mult_2.MULT_BYPASS = "DISABLED";
    defparam mult_11_mult_2.RESETMODE = "SYNC";
    CCU2C rem_10_add_1311_15 (.A0(n13600), .B0(n28359), .C0(n1907[28]), 
          .D0(n38291), .A1(n13600), .B1(n28359), .C1(n1907[29]), .D1(n38290), 
          .CIN(n30596), .COUT(n30597), .S0(n2006[28]), .S1(n2006[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1311_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1311_15.INJECT1_0 = "NO";
    defparam rem_10_add_1311_15.INJECT1_1 = "NO";
    LUT4 rem_10_i2261_3_lut (.A(n3336), .B(n3392_adj_2163[21]), .C(n3359), 
         .Z(n3435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2261_3_lut.init = 16'hcaca;
    CCU2C div_9_add_1512_7 (.A0(n13590), .B0(n28440), .C0(n2204[18]), 
          .D0(n2151), .A1(n13590), .B1(n28440), .C1(n2204[19]), .D1(n2150), 
          .CIN(n30682), .COUT(n30683), .S0(n2303[18]), .S1(n2303[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1512_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1512_7.INJECT1_0 = "NO";
    defparam div_9_add_1512_7.INJECT1_1 = "NO";
    CCU2C div_9_add_2182_9 (.A0(n13547), .B0(n28588), .C0(n3194[10]), 
          .D0(n3149), .A1(n13547), .B1(n28588), .C1(n3194[11]), .D1(n3148), 
          .CIN(n30803), .COUT(n30804), .S0(n3293[10]), .S1(n3293[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_9.INIT0 = 16'hf1e0;
    defparam div_9_add_2182_9.INIT1 = 16'hf1e0;
    defparam div_9_add_2182_9.INJECT1_0 = "NO";
    defparam div_9_add_2182_9.INJECT1_1 = "NO";
    LUT4 rem_10_i2263_3_lut (.A(n3338), .B(n3392_adj_2163[19]), .C(n3359), 
         .Z(n3437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2263_3_lut.init = 16'hcaca;
    CCU2C rem_10_add_1311_13 (.A0(n13600), .B0(n28359), .C0(n1907[26]), 
          .D0(n1846), .A1(n13600), .B1(n28359), .C1(n1907[27]), .D1(n1845), 
          .CIN(n30595), .COUT(n30596), .S0(n2006[26]), .S1(n2006[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1311_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1311_13.INJECT1_0 = "NO";
    defparam rem_10_add_1311_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1922_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[25]), 
         .D(n38235), .Z(n2936)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1922_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2269_3_lut (.A(n3344), .B(n3392_adj_2163[13]), .C(n3359), 
         .Z(n3443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2269_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1918_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[29]), 
         .D(n2833), .Z(n2932)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1918_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_26227_11 (.A0(n13629), .B0(n28492), .C0(n3293[11]), .D0(n3247), 
          .A1(n13629), .B1(n28492), .C1(n3293[12]), .D1(n3246_adj_548), 
          .CIN(n30537), .COUT(n30538), .S0(n3392[11]), .S1(n3392[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_11.INIT0 = 16'h0e1f;
    defparam add_26227_11.INIT1 = 16'h0e1f;
    defparam add_26227_11.INJECT1_0 = "NO";
    defparam add_26227_11.INJECT1_1 = "NO";
    LUT4 rem_10_i2201_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[14]), 
         .D(n3244_adj_551), .Z(n3343)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2201_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1311_11 (.A0(n13600), .B0(n28359), .C0(n1907[24]), 
          .D0(n1848), .A1(n13600), .B1(n28359), .C1(n1907[25]), .D1(n1847), 
          .CIN(n30594), .COUT(n30595), .S0(n2006[24]), .S1(n2006[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_11.INIT0 = 16'hf1e0;
    defparam rem_10_add_1311_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1311_11.INJECT1_0 = "NO";
    defparam rem_10_add_1311_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1512_5 (.A0(n13590), .B0(n28440), .C0(n2204[16]), 
          .D0(n2153), .A1(n13590), .B1(n28440), .C1(n2204[17]), .D1(n38278), 
          .CIN(n30681), .COUT(n30682), .S0(n2303[16]), .S1(n2303[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1512_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1512_5.INJECT1_0 = "NO";
    defparam div_9_add_1512_5.INJECT1_1 = "NO";
    CCU2C add_26227_9 (.A0(n13629), .B0(n28492), .C0(n3293[9]), .D0(n3249), 
          .A1(n13629), .B1(n28492), .C1(n3293[10]), .D1(n3248), .CIN(n30536), 
          .COUT(n30537), .S0(n3392[9]), .S1(n3392[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_9.INIT0 = 16'hf1e0;
    defparam add_26227_9.INIT1 = 16'hf1e0;
    defparam add_26227_9.INJECT1_0 = "NO";
    defparam add_26227_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1311_9 (.A0(n13600), .B0(n28359), .C0(n1907[22]), 
          .D0(n1850), .A1(n13600), .B1(n28359), .C1(n1907[23]), .D1(n1849), 
          .CIN(n30593), .COUT(n30594), .S0(n2006[22]), .S1(n2006[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1311_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1311_9.INJECT1_0 = "NO";
    defparam rem_10_add_1311_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1311_7 (.A0(n13600), .B0(n28359), .C0(n1907[20]), 
          .D0(n38292), .A1(n13600), .B1(n28359), .C1(n1907[21]), .D1(n1851), 
          .CIN(n30592), .COUT(n30593), .S0(n2006[20]), .S1(n2006[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_7.INIT0 = 16'hf1e0;
    defparam rem_10_add_1311_7.INIT1 = 16'h0e1f;
    defparam rem_10_add_1311_7.INJECT1_0 = "NO";
    defparam rem_10_add_1311_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1512_3 (.A0(n13590), .B0(n28440), .C0(n2204[14]), 
          .D0(n337), .A1(n13590), .B1(n28440), .C1(n2204[15]), .D1(n2154), 
          .CIN(n30680), .COUT(n30681), .S0(n2303[14]), .S1(n2303[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1512_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1512_3.INJECT1_0 = "NO";
    defparam div_9_add_1512_3.INJECT1_1 = "NO";
    CCU2C div_9_add_2182_7 (.A0(n13547), .B0(n28588), .C0(n3194[8]), .D0(n38202), 
          .A1(n13547), .B1(n28588), .C1(n3194[9]), .D1(n3150), .CIN(n30802), 
          .COUT(n30803), .S0(n3293[8]), .S1(n3293[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_7.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_7.INIT1 = 16'hf1e0;
    defparam div_9_add_2182_7.INJECT1_0 = "NO";
    defparam div_9_add_2182_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1847_5 (.A0(n13624), .B0(n28462), .C0(n2699[11]), 
          .D0(n2653), .A1(n13624), .B1(n28462), .C1(n2699[12]), .D1(n2652), 
          .CIN(n30974), .COUT(n30975), .S0(n2798[11]), .S1(n2798[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1847_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1847_5.INJECT1_0 = "NO";
    defparam div_13_add_1847_5.INJECT1_1 = "NO";
    CCU2C add_26227_7 (.A0(n13629), .B0(n28492), .C0(n3293[7]), .D0(n38196), 
          .A1(n13629), .B1(n28492), .C1(n3293[8]), .D1(n3250_adj_554), 
          .CIN(n30535), .COUT(n30536), .S0(n3392[7]), .S1(n3392[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_7.INIT0 = 16'h0e1f;
    defparam add_26227_7.INIT1 = 16'hf1e0;
    defparam add_26227_7.INJECT1_0 = "NO";
    defparam add_26227_7.INJECT1_1 = "NO";
    LUT4 rem_10_i1931_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[16]), 
         .D(n2846), .Z(n2945)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1931_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1940_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[7]), 
         .D(n593), .Z(n2954)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1940_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2266_3_lut (.A(n3341), .B(n3392_adj_2163[16]), .C(n3359), 
         .Z(n3440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2266_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2262_3_lut (.A(n3337), .B(n3392_adj_2163[20]), .C(n3359), 
         .Z(n3436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2262_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2267_3_lut (.A(n3342), .B(n3392_adj_2163[15]), .C(n3359), 
         .Z(n3441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2267_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1937_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[10]), 
         .D(n38237), .Z(n2951)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1937_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1847_3 (.A0(n13624), .B0(n28462), .C0(n2699[9]), 
          .D0(n342), .A1(n13624), .B1(n28462), .C1(n2699[10]), .D1(n2654), 
          .CIN(n30973), .COUT(n30974), .S0(n2798[9]), .S1(n2798[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1847_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_3.INJECT1_0 = "NO";
    defparam div_13_add_1847_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_16 (.A(n38179), .B(n38175), .C(n3449), .D(n3447), 
         .Z(n33580)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_16.init = 16'h8000;
    CCU2C add_26227_5 (.A0(n13629), .B0(n28492), .C0(n3293[5]), .D0(n3253), 
          .A1(n13629), .B1(n28492), .C1(n3293[6]), .D1(n3252), .CIN(n30534), 
          .COUT(n30535), .S0(n3392[5]), .S1(n3392[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_5.INIT0 = 16'hf1e0;
    defparam add_26227_5.INIT1 = 16'hf1e0;
    defparam add_26227_5.INJECT1_0 = "NO";
    defparam add_26227_5.INJECT1_1 = "NO";
    LUT4 rem_10_i2197_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[18]), 
         .D(n3240_adj_561), .Z(n3339)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2197_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_17 (.A(n34976), .B(n38059), .C(n3428), .D(n3444), 
         .Z(n39_adj_523)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_17.init = 16'hfffe;
    LUT4 i1_4_lut_adj_18 (.A(n38186), .B(n3425), .C(n3392_adj_2163[26]), 
         .D(n3359), .Z(n34976)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_18.init = 16'hfcee;
    LUT4 div_13_i2197_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[18]), 
         .D(n3240_adj_564), .Z(n3339_adj_565)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2197_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2254_3_lut (.A(n38184), .B(n3392_adj_2163[28]), .C(n3359), 
         .Z(n3428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2254_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2193_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[22]), 
         .D(n3236_adj_568), .Z(n3335)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2193_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1933_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[14]), 
         .D(n2848_adj_570), .Z(n2947_adj_571)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1933_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2270_3_lut (.A(n3345), .B(n3392_adj_2163[12]), .C(n3359), 
         .Z(n3444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2270_3_lut.init = 16'hcaca;
    CCU2C add_26227_3 (.A0(n13629), .B0(n28492), .C0(n3293[3]), .D0(n348), 
          .A1(n13629), .B1(n28492), .C1(n3293[4]), .D1(n3254), .CIN(n30533), 
          .COUT(n30534), .S0(n3392[3]), .S1(n3392[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_3.INIT0 = 16'hf1e0;
    defparam add_26227_3.INIT1 = 16'h0e1f;
    defparam add_26227_3.INJECT1_0 = "NO";
    defparam add_26227_3.INJECT1_1 = "NO";
    CCU2C add_26227_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n12154), .B1(n5), .C1(distance[0]), .D1(n35[2]), .COUT(n30533));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_26227_1.INIT0 = 16'h0000;
    defparam add_26227_1.INIT1 = 16'habef;
    defparam add_26227_1.INJECT1_0 = "NO";
    defparam add_26227_1.INJECT1_1 = "NO";
    LUT4 rem_10_i2251_3_lut (.A(n3326), .B(n3392_adj_2163[31]), .C(n3359), 
         .Z(n3425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2251_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1934_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[13]), 
         .D(n2849), .Z(n2948)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1934_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_842_Select_2_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[2]), 
         .D(n2983), .Z(duty0_14__N_410[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_2_i4_3_lut_4_lut.init = 16'hff10;
    LUT4 select_842_Select_1_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[1]), 
         .D(n2983), .Z(duty0_14__N_410[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_1_i4_3_lut_4_lut.init = 16'hff10;
    LUT4 i22780_2_lut_4_lut (.A(n1), .B(n13790), .C(n89[0]), .D(n197[8]), 
         .Z(duty3_14__N_488[8])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i22780_2_lut_4_lut.init = 16'h2000;
    CCU2C div_9_add_2182_5 (.A0(n13547), .B0(n28588), .C0(n3194[6]), .D0(n3153), 
          .A1(n13547), .B1(n28588), .C1(n3194[7]), .D1(n3152), .CIN(n30801), 
          .COUT(n30802), .S0(n3293[6]), .S1(n3293[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_5.INIT0 = 16'hf1e0;
    defparam div_9_add_2182_5.INIT1 = 16'hf1e0;
    defparam div_9_add_2182_5.INJECT1_0 = "NO";
    defparam div_9_add_2182_5.INJECT1_1 = "NO";
    LUT4 rem_10_i2273_3_lut (.A(n3348), .B(n3392_adj_2163[9]), .C(n3359), 
         .Z(n3447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2273_3_lut.init = 16'hcaca;
    CCU2C div_9_add_1512_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n51), .D1(n35[13]), 
          .COUT(n30680), .S1(n2303[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1512_1.INIT0 = 16'h0000;
    defparam div_9_add_1512_1.INIT1 = 16'habef;
    defparam div_9_add_1512_1.INJECT1_0 = "NO";
    defparam div_9_add_1512_1.INJECT1_1 = "NO";
    LUT4 rem_10_i2186_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[29]), 
         .D(n3229), .Z(n3328)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2186_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1935_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[12]), 
         .D(n2850), .Z(n2949)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1935_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2200_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[15]), 
         .D(n3243_adj_580), .Z(n3342)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2200_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2343_3_lut (.A(n3450), .B(n38178), .C(n3458), .Z(n3549)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2343_3_lut.init = 16'h9a9a;
    LUT4 rem_10_i1936_3_lut_4_lut (.A(n28307), .B(n13598), .C(n2897_adj_2162[11]), 
         .D(n2851), .Z(n2950)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1936_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_19 (.A(n36114), .B(n36120), .C(n36110), .D(n36116), 
         .Z(n13629)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_19.init = 16'hfffe;
    LUT4 i1_4_lut_adj_20 (.A(n3235), .B(n3241_adj_532), .C(n3242), .D(n3231), 
         .Z(n36114)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_20.init = 16'hfffe;
    LUT4 i1_4_lut_adj_21 (.A(n3232), .B(n36112), .C(n36090), .D(n3240), 
         .Z(n36120)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_21.init = 16'hfffe;
    LUT4 i1_4_lut_adj_22 (.A(n3243), .B(n3233_adj_522), .C(n3246_adj_548), 
         .D(n3227), .Z(n36110)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_22.init = 16'hfffe;
    LUT4 i1_4_lut_adj_23 (.A(n3244), .B(n3245), .C(n3236), .D(n3230), 
         .Z(n36116)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_23.init = 16'hfffe;
    LUT4 rem_10_i2344_4_lut (.A(n3451), .B(n3452), .C(n3458), .D(n3453), 
         .Z(n3550)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2344_4_lut.init = 16'h6aaa;
    LUT4 i1_4_lut_adj_24 (.A(n3237), .B(n3239), .C(n3228), .D(n3238), 
         .Z(n36112)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_24.init = 16'hfffe;
    LUT4 rem_10_i2345_3_lut (.A(n3452), .B(n3453), .C(n3458), .Z(n3551)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2345_3_lut.init = 16'h6a6a;
    LUT4 i1_4_lut_adj_25 (.A(n35824), .B(n35786), .C(n3250_adj_554), .D(n28176), 
         .Z(n28492)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_25.init = 16'ha8a0;
    LUT4 rem_10_i2339_3_lut (.A(n3446), .B(n33580), .C(n3458), .Z(n3545)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2339_3_lut.init = 16'h9a9a;
    LUT4 i1_3_lut_adj_26 (.A(n3247), .B(n3248), .C(n3249), .Z(n35824)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_26.init = 16'h8080;
    LUT4 rem_10_i2280_3_lut (.A(n598), .B(n3392_adj_2163[2]), .C(n3359), 
         .Z(n3454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2280_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2185_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[30]), 
         .D(n3228_adj_582), .Z(n3327)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24224_3_lut (.A(n348), .B(n3253), .C(n3254), .Z(n28176)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24224_3_lut.init = 16'hecec;
    LUT4 i1_3_lut_adj_27 (.A(n27382), .B(n3), .C(n48), .Z(duty0_14__N_426[12])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_27.init = 16'h2020;
    LUT4 i1_4_lut_adj_28 (.A(n2039), .B(n34486), .C(n36046), .D(n2042), 
         .Z(n13605)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_28.init = 16'hfffe;
    LUT4 rem_10_i2184_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[31]), 
         .D(n3227_adj_584), .Z(n3326)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_29 (.A(n2045), .B(n2043), .C(n2044), .D(n2041), 
         .Z(n34486)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_29.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_30 (.A(n38232), .B(n2798[18]), .C(n38228), 
         .D(n2845_adj_585), .Z(n35452)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_30.init = 16'hffca;
    CCU2C div_9_add_2182_3 (.A0(n13547), .B0(n28588), .C0(n3194[4]), .D0(n347), 
          .A1(n13547), .B1(n28588), .C1(n3194[5]), .D1(n3154), .CIN(n30800), 
          .COUT(n30801), .S0(n3293[4]), .S1(n3293[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_3.INIT0 = 16'hf1e0;
    defparam div_9_add_2182_3.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_3.INJECT1_0 = "NO";
    defparam div_9_add_2182_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1847_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n343), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30973), .S1(n2798[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_1.INIT0 = 16'h0000;
    defparam div_13_add_1847_1.INIT1 = 16'h555a;
    defparam div_13_add_1847_1.INJECT1_0 = "NO";
    defparam div_13_add_1847_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1445_19 (.A0(n13605), .B0(n28263), .C0(n2105[31]), 
          .D0(n2039), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30679), .S0(n2204[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1445_19.INIT1 = 16'h0000;
    defparam div_9_add_1445_19.INJECT1_0 = "NO";
    defparam div_9_add_1445_19.INJECT1_1 = "NO";
    LUT4 i24524_2_lut_rep_223 (.A(n28468), .B(n13622), .Z(n38228)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24524_2_lut_rep_223.init = 16'heeee;
    LUT4 i1_4_lut_adj_31 (.A(n2047), .B(n28247), .C(n2048), .D(n2049), 
         .Z(n28263)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_31.init = 16'h8000;
    CCU2C div_13_add_1780_23 (.A0(n13625), .B0(n28456), .C0(n2600[30]), 
          .D0(n2535), .A1(n13625), .B1(n28456), .C1(n2600[31]), .D1(n2534), 
          .CIN(n30971), .S0(n2699[30]), .S1(n2699[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_23.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_23.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_23.INJECT1_0 = "NO";
    defparam div_13_add_1780_23.INJECT1_1 = "NO";
    LUT4 rem_10_i2209_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[6]), 
         .D(n38198), .Z(n3351)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2209_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1780_21 (.A0(n13625), .B0(n28456), .C0(n2600[28]), 
          .D0(n2537), .A1(n13625), .B1(n28456), .C1(n2600[29]), .D1(n2536), 
          .CIN(n30970), .COUT(n30971), .S0(n2699[28]), .S1(n2699[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_21.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_21.INJECT1_0 = "NO";
    defparam div_13_add_1780_21.INJECT1_1 = "NO";
    LUT4 i24294_4_lut (.A(n2051), .B(n2050), .C(n27986), .D(n2052), 
         .Z(n28247)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24294_4_lut.init = 16'heccc;
    LUT4 div_13_i1862_3_lut_rep_222_4_lut (.A(n28468), .B(n13622), .C(n2798[18]), 
         .D(n38232), .Z(n38227)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1862_3_lut_rep_222_4_lut.init = 16'hf1e0;
    LUT4 i24036_3_lut (.A(n336), .B(n2053), .C(n2054), .Z(n27986)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24036_3_lut.init = 16'hecec;
    LUT4 rem_10_i2199_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[16]), 
         .D(n3242_adj_588), .Z(n3341)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2199_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2182_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[3]), .D1(duty0_14__N_426[1]), 
          .COUT(n30800), .S1(n3293[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_1.INIT0 = 16'h0000;
    defparam div_9_add_2182_1.INIT1 = 16'h04bf;
    defparam div_9_add_2182_1.INJECT1_0 = "NO";
    defparam div_9_add_2182_1.INJECT1_1 = "NO";
    LUT4 div_13_i1856_3_lut_rep_217_4_lut (.A(n28468), .B(n13622), .C(n2798[24]), 
         .D(n2739), .Z(n38222)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1856_3_lut_rep_217_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1780_19 (.A0(n13625), .B0(n28456), .C0(n2600[26]), 
          .D0(n2539), .A1(n13625), .B1(n28456), .C1(n2600[27]), .D1(n2538), 
          .CIN(n30969), .COUT(n30970), .S0(n2699[26]), .S1(n2699[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_19.INJECT1_0 = "NO";
    defparam div_13_add_1780_19.INJECT1_1 = "NO";
    PFUMX pwm_cnt_14__I_0_51_i24 (.BLUT(n16_adj_589), .ALUT(n22), .C0(n36923), 
          .Z(n24)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    CCU2C rem_10_add_1311_5 (.A0(n13600), .B0(n28359), .C0(n1907[18]), 
          .D0(n1854), .A1(n13600), .B1(n28359), .C1(n1907[19]), .D1(n1853), 
          .CIN(n30591), .COUT(n30592), .S0(n2006[18]), .S1(n2006[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_5.INIT0 = 16'h0e1f;
    defparam rem_10_add_1311_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1311_5.INJECT1_0 = "NO";
    defparam rem_10_add_1311_5.INJECT1_1 = "NO";
    CCU2C add_26228_29 (.A0(n3556), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n3556), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30528), 
          .S0(n38[27]), .S1(n38[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_29.INIT0 = 16'h5550;
    defparam add_26228_29.INIT1 = 16'h5550;
    defparam add_26228_29.INJECT1_0 = "NO";
    defparam add_26228_29.INJECT1_1 = "NO";
    LUT4 div_13_i1871_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[9]), 
         .D(n2754), .Z(n2853_adj_591)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1871_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1780_17 (.A0(n13625), .B0(n28456), .C0(n2600[24]), 
          .D0(n2541), .A1(n13625), .B1(n28456), .C1(n2600[25]), .D1(n2540), 
          .CIN(n30968), .COUT(n30969), .S0(n2699[24]), .S1(n2699[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_17.INJECT1_0 = "NO";
    defparam div_13_add_1780_17.INJECT1_1 = "NO";
    LUT4 div_13_i1858_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[22]), 
         .D(n2741), .Z(n2840)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1858_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1850_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[30]), 
         .D(n2733), .Z(n2832_adj_592)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1850_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1445_17 (.A0(n13605), .B0(n28263), .C0(n2105[29]), 
          .D0(n2041), .A1(n13605), .B1(n28263), .C1(n2105[30]), .D1(n2040), 
          .CIN(n30678), .COUT(n30679), .S0(n2204[29]), .S1(n2204[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1445_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1445_17.INJECT1_0 = "NO";
    defparam div_9_add_1445_17.INJECT1_1 = "NO";
    CCU2C div_9_add_1445_15 (.A0(n13605), .B0(n28263), .C0(n2105[27]), 
          .D0(n2043), .A1(n13605), .B1(n28263), .C1(n2105[28]), .D1(n2042), 
          .CIN(n30677), .COUT(n30678), .S0(n2204[27]), .S1(n2204[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1445_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1445_15.INJECT1_0 = "NO";
    defparam div_9_add_1445_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_1311_3 (.A0(n12154), .B0(n5), .C0(n42), .D0(n2[16]), 
          .A1(n13600), .B1(n28359), .C1(n1907[17]), .D1(n583), .CIN(n30590), 
          .COUT(n30591), .S0(n2006[16]), .S1(n2006[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_3.INIT0 = 16'h5410;
    defparam rem_10_add_1311_3.INIT1 = 16'hf1e0;
    defparam rem_10_add_1311_3.INJECT1_0 = "NO";
    defparam rem_10_add_1311_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1780_15 (.A0(n13625), .B0(n28456), .C0(n2600[22]), 
          .D0(n2543), .A1(n13625), .B1(n28456), .C1(n2600[23]), .D1(n2542), 
          .CIN(n30967), .COUT(n30968), .S0(n2699[22]), .S1(n2699[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_15.INJECT1_0 = "NO";
    defparam div_13_add_1780_15.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_29 (.A0(n13548), .B0(n28578), .C0(n3095[31]), 
          .D0(n3029), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30799), .S0(n3194[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_29.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_29.INIT1 = 16'h0000;
    defparam div_9_add_2115_29.INJECT1_0 = "NO";
    defparam div_9_add_2115_29.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_32 (.A(n27382), .B(n3), .C(n75_adj_1), .Z(duty0_14__N_426[3])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_32.init = 16'h2020;
    CCU2C div_9_add_2115_27 (.A0(n13548), .B0(n28578), .C0(n3095[29]), 
          .D0(n38211), .A1(n13548), .B1(n28578), .C1(n3095[30]), .D1(n38212), 
          .CIN(n30798), .COUT(n30799), .S0(n3194[29]), .S1(n3194[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_27.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_27.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_27.INJECT1_0 = "NO";
    defparam div_9_add_2115_27.INJECT1_1 = "NO";
    CCU2C rem_10_add_1311_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n45), .D1(n2[15]), 
          .COUT(n30590));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1311_1.INIT0 = 16'h000F;
    defparam rem_10_add_1311_1.INIT1 = 16'habef;
    defparam rem_10_add_1311_1.INJECT1_0 = "NO";
    defparam rem_10_add_1311_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_33 (.A(n35684), .B(n35678), .C(n2545), .D(n2542), 
         .Z(n13625)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_33.init = 16'hfffe;
    LUT4 i1_4_lut_adj_34 (.A(n2541), .B(n35680), .C(n2543), .D(n2536), 
         .Z(n35684)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_34.init = 16'hfffe;
    CCU2C add_26228_27 (.A0(n66_adj_2), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n63_adj_3), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30527), .COUT(n30528), .S0(n38[25]), .S1(n38[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_27.INIT0 = 16'h5550;
    defparam add_26228_27.INIT1 = 16'h5550;
    defparam add_26228_27.INJECT1_0 = "NO";
    defparam add_26228_27.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_35 (.A(n2540), .B(n2535), .C(n2544), .D(n2539), 
         .Z(n35678)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_35.init = 16'hfffe;
    LUT4 div_13_i1863_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[17]), 
         .D(n2746), .Z(n2845_adj_585)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1863_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2211_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[4]), 
         .D(n3254_adj_597), .Z(n3353)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2211_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2115_25 (.A0(n13548), .B0(n28578), .C0(n3095[27]), 
          .D0(n3033), .A1(n13548), .B1(n28578), .C1(n3095[28]), .D1(n3032), 
          .CIN(n30797), .COUT(n30798), .S0(n3194[27]), .S1(n3194[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_25.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_25.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_25.INJECT1_0 = "NO";
    defparam div_9_add_2115_25.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_23 (.A0(n13548), .B0(n28578), .C0(n3095[25]), 
          .D0(n3035), .A1(n13548), .B1(n28578), .C1(n3095[26]), .D1(n3034), 
          .CIN(n30796), .COUT(n30797), .S0(n3194[25]), .S1(n3194[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_23.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_23.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_23.INJECT1_0 = "NO";
    defparam div_9_add_2115_23.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_36 (.A(n2538), .B(n2534), .C(n2546), .D(n2537), 
         .Z(n35680)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_36.init = 16'hfffe;
    LUT4 rem_10_i2204_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[11]), 
         .D(n3247_adj_599), .Z(n3346)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2204_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23478_2_lut_rep_311 (.A(n60_adj_4), .B(n3), .Z(n38316)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23478_2_lut_rep_311.init = 16'heeee;
    LUT4 div_13_i1872_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[8]), 
         .D(n343), .Z(n2854_adj_601)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1872_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1445_13 (.A0(n13605), .B0(n28263), .C0(n2105[25]), 
          .D0(n2045), .A1(n13605), .B1(n28263), .C1(n2105[26]), .D1(n2044), 
          .CIN(n30676), .COUT(n30677), .S0(n2204[25]), .S1(n2204[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1445_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1445_13.INJECT1_0 = "NO";
    defparam div_9_add_1445_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1780_13 (.A0(n13625), .B0(n28456), .C0(n2600[20]), 
          .D0(n2545), .A1(n13625), .B1(n28456), .C1(n2600[21]), .D1(n2544), 
          .CIN(n30966), .COUT(n30967), .S0(n2699[20]), .S1(n2699[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_13.INJECT1_0 = "NO";
    defparam div_13_add_1780_13.INJECT1_1 = "NO";
    LUT4 i23441_2_lut_3_lut (.A(n60_adj_4), .B(n3), .C(n27382), .Z(duty0_14__N_426[8])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23441_2_lut_3_lut.init = 16'he0e0;
    LUT4 i23475_2_lut_rep_312 (.A(n57), .B(n3), .Z(n38317)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23475_2_lut_rep_312.init = 16'heeee;
    LUT4 i23440_2_lut_3_lut (.A(n57), .B(n3), .C(n27382), .Z(duty0_14__N_426[9])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23440_2_lut_3_lut.init = 16'he0e0;
    CCU2C div_9_add_2115_21 (.A0(n13548), .B0(n28578), .C0(n3095[23]), 
          .D0(n3037), .A1(n13548), .B1(n28578), .C1(n3095[24]), .D1(n3036), 
          .CIN(n30795), .COUT(n30796), .S0(n3194[23]), .S1(n3194[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_21.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_21.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_21.INJECT1_0 = "NO";
    defparam div_9_add_2115_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_37 (.A(n2548), .B(n28299), .C(n2547), .D(n2549), 
         .Z(n28456)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_37.init = 16'h8000;
    LUT4 div_13_i2199_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[16]), 
         .D(n3242_adj_603), .Z(n3341_adj_604)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2199_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24346_4_lut (.A(n2551), .B(n2550), .C(n28048), .D(n2552), 
         .Z(n28299)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24346_4_lut.init = 16'heccc;
    CCU2C div_9_add_2115_19 (.A0(n13548), .B0(n28578), .C0(n3095[21]), 
          .D0(n3039), .A1(n13548), .B1(n28578), .C1(n3095[22]), .D1(n3038), 
          .CIN(n30794), .COUT(n30795), .S0(n3194[21]), .S1(n3194[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_19.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_19.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_19.INJECT1_0 = "NO";
    defparam div_9_add_2115_19.INJECT1_1 = "NO";
    LUT4 i24098_3_lut (.A(n341_adj_605), .B(n2553), .C(n2554), .Z(n28048)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24098_3_lut.init = 16'hecec;
    CCU2C div_13_add_1780_11 (.A0(n13625), .B0(n28456), .C0(n2600[18]), 
          .D0(n2547), .A1(n13625), .B1(n28456), .C1(n2600[19]), .D1(n2546), 
          .CIN(n30965), .COUT(n30966), .S0(n2699[18]), .S1(n2699[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_11.INJECT1_0 = "NO";
    defparam div_13_add_1780_11.INJECT1_1 = "NO";
    LUT4 rem_10_i2208_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[7]), 
         .D(n3251), .Z(n3350)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2208_3_lut_4_lut.init = 16'hf1e0;
    PFUMX pwm_cnt_14__I_0_52_i24 (.BLUT(n16_adj_607), .ALUT(n22_adj_608), 
          .C0(n36866), .Z(n24_adj_609)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    LUT4 div_13_i1865_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[15]), 
         .D(n2748), .Z(n2847_adj_610)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1865_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1851_3_lut_rep_214_4_lut (.A(n28468), .B(n13622), .C(n2798[29]), 
         .D(n2734), .Z(n38219)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1851_3_lut_rep_214_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1445_11 (.A0(n13605), .B0(n28263), .C0(n2105[23]), 
          .D0(n2047), .A1(n13605), .B1(n28263), .C1(n2105[24]), .D1(n38281), 
          .CIN(n30675), .COUT(n30676), .S0(n2204[23]), .S1(n2204[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1445_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1445_11.INJECT1_0 = "NO";
    defparam div_9_add_1445_11.INJECT1_1 = "NO";
    LUT4 div_13_i2188_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[27]), 
         .D(n3231_adj_612), .Z(n3330_adj_613)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2212_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[3]), 
         .D(n597), .Z(n3354)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2212_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1849_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[31]), 
         .D(n2732), .Z(n2831)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1849_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1864_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[16]), 
         .D(n2747), .Z(n2846_adj_615)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1864_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1780_9 (.A0(n13625), .B0(n28456), .C0(n2600[16]), 
          .D0(n2549), .A1(n13625), .B1(n28456), .C1(n2600[17]), .D1(n2548), 
          .CIN(n30964), .COUT(n30965), .S0(n2699[16]), .S1(n2699[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1780_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1780_9.INJECT1_0 = "NO";
    defparam div_13_add_1780_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1780_7 (.A0(n13625), .B0(n28456), .C0(n2600[14]), 
          .D0(n2551), .A1(n13625), .B1(n28456), .C1(n2600[15]), .D1(n2550), 
          .CIN(n30963), .COUT(n30964), .S0(n2699[14]), .S1(n2699[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1780_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1780_7.INJECT1_0 = "NO";
    defparam div_13_add_1780_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1445_9 (.A0(n13605), .B0(n28263), .C0(n2105[21]), 
          .D0(n2049), .A1(n13605), .B1(n28263), .C1(n2105[22]), .D1(n2048), 
          .CIN(n30674), .COUT(n30675), .S0(n2204[21]), .S1(n2204[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1445_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1445_9.INJECT1_0 = "NO";
    defparam div_9_add_1445_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1780_5 (.A0(n13625), .B0(n28456), .C0(n2600[12]), 
          .D0(n2553), .A1(n13625), .B1(n28456), .C1(n2600[13]), .D1(n2552), 
          .CIN(n30962), .COUT(n30963), .S0(n2699[12]), .S1(n2699[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1780_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1780_5.INJECT1_0 = "NO";
    defparam div_13_add_1780_5.INJECT1_1 = "NO";
    CCU2C div_13_add_1780_3 (.A0(n13625), .B0(n28456), .C0(n2600[10]), 
          .D0(n341_adj_605), .A1(n13625), .B1(n28456), .C1(n2600[11]), 
          .D1(n2554), .CIN(n30961), .COUT(n30962), .S0(n2699[10]), .S1(n2699[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1780_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1780_3.INJECT1_0 = "NO";
    defparam div_13_add_1780_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1780_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n342), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30961), .S1(n2699[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1780_1.INIT0 = 16'h0000;
    defparam div_13_add_1780_1.INIT1 = 16'h555a;
    defparam div_13_add_1780_1.INJECT1_0 = "NO";
    defparam div_13_add_1780_1.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_17 (.A0(n13548), .B0(n28578), .C0(n3095[19]), 
          .D0(n3041), .A1(n13548), .B1(n28578), .C1(n3095[20]), .D1(n3040), 
          .CIN(n30793), .COUT(n30794), .S0(n3194[19]), .S1(n3194[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_17.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_17.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_17.INJECT1_0 = "NO";
    defparam div_9_add_2115_17.INJECT1_1 = "NO";
    LUT4 div_13_i1859_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[21]), 
         .D(n2742), .Z(n2841_adj_616)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1859_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2205_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[10]), 
         .D(n3248_adj_618), .Z(n3347)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2205_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1870_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[10]), 
         .D(n2753), .Z(n2852)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1870_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1713_23 (.A0(n13627), .B0(n28446), .C0(n2501[31]), 
          .D0(n38254), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30960), .S0(n2600[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_23.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_23.INIT1 = 16'h0000;
    defparam div_13_add_1713_23.INJECT1_0 = "NO";
    defparam div_13_add_1713_23.INJECT1_1 = "NO";
    LUT4 div_13_i1853_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[27]), 
         .D(n2736), .Z(n2835_adj_619)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1853_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1860_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[20]), 
         .D(n2743), .Z(n2842_adj_620)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1860_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2206_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[9]), 
         .D(n3249_adj_622), .Z(n3348)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2206_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2115_15 (.A0(n13548), .B0(n28578), .C0(n3095[17]), 
          .D0(n3043), .A1(n13548), .B1(n28578), .C1(n3095[18]), .D1(n3042), 
          .CIN(n30792), .COUT(n30793), .S0(n3194[17]), .S1(n3194[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_15.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_15.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_15.INJECT1_0 = "NO";
    defparam div_9_add_2115_15.INJECT1_1 = "NO";
    LUT4 rem_10_i2196_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[19]), 
         .D(n3239_adj_624), .Z(n3338)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2196_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1713_21 (.A0(n13627), .B0(n28446), .C0(n2501[29]), 
          .D0(n2437), .A1(n13627), .B1(n28446), .C1(n2501[30]), .D1(n2436), 
          .CIN(n30959), .COUT(n30960), .S0(n2600[29]), .S1(n2600[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_21.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_21.INJECT1_0 = "NO";
    defparam div_13_add_1713_21.INJECT1_1 = "NO";
    PFUMX pwm_cnt_14__I_0_53_i24 (.BLUT(n16_adj_625), .ALUT(n22_adj_626), 
          .C0(n36809), .Z(n24_adj_627)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    CCU2C div_9_add_1445_7 (.A0(n13605), .B0(n28263), .C0(n2105[19]), 
          .D0(n2051), .A1(n13605), .B1(n28263), .C1(n2105[20]), .D1(n2050), 
          .CIN(n30673), .COUT(n30674), .S0(n2204[19]), .S1(n2204[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1445_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1445_7.INJECT1_0 = "NO";
    defparam div_9_add_1445_7.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_13 (.A0(n13548), .B0(n28578), .C0(n3095[15]), 
          .D0(n3045), .A1(n13548), .B1(n28578), .C1(n3095[16]), .D1(n3044), 
          .CIN(n30791), .COUT(n30792), .S0(n3194[15]), .S1(n3194[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_13.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_13.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_13.INJECT1_0 = "NO";
    defparam div_9_add_2115_13.INJECT1_1 = "NO";
    LUT4 div_13_i1854_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[26]), 
         .D(n2737), .Z(n2836_adj_628)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1854_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2191_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[24]), 
         .D(n3234_adj_630), .Z(n3333)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1867_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[13]), 
         .D(n2750), .Z(n2849_adj_631)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1867_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3399_bdd_4_lut (.A(n3327_adj_632), .B(n3332_adj_633), .C(n3345_adj_634), 
         .D(n3335_adj_635), .Z(n37516)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3399_bdd_4_lut.init = 16'hfffe;
    LUT4 div_13_i1868_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[12]), 
         .D(n2751), .Z(n2850_adj_636)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1868_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1861_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[19]), 
         .D(n2744), .Z(n2843_adj_637)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1861_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2195_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[20]), 
         .D(n3238_adj_639), .Z(n3337)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2195_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32216_4_lut (.A(n38398), .B(n38397), .C(n38396), .D(n36909), 
         .Z(n36923)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32216_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_38 (.A(n36010), .B(n36000), .C(n3036), .D(n3041), 
         .Z(n13548)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_38.init = 16'hfffe;
    LUT4 div_13_i2411_3_lut_4_lut (.A(n28468), .B(n13622), .C(n3556), 
         .D(n4990[7]), .Z(n197[7])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2411_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i1_4_lut_adj_39 (.A(n36008), .B(n3043), .C(n35982), .D(n3045), 
         .Z(n36010)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_39.init = 16'hfffe;
    LUT4 i1_4_lut_adj_40 (.A(n3034), .B(n3032), .C(n3042), .D(n3046), 
         .Z(n36000)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_40.init = 16'hfffe;
    LUT4 i1_4_lut_adj_41 (.A(n35992), .B(n36002), .C(n3029), .D(n3037), 
         .Z(n36008)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_41.init = 16'hfffe;
    LUT4 div_13_i1852_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[28]), 
         .D(n2735), .Z(n2834_adj_640)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1852_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2202_3_lut_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[13]), 
         .D(n3245_adj_642), .Z(n3344)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2202_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1857_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[23]), 
         .D(n38233), .Z(n2839_adj_643)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1857_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1855_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[25]), 
         .D(n2738), .Z(n2837)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1855_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_42 (.A(n3033), .B(n3038), .C(n3044), .D(n3040), 
         .Z(n36002)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_42.init = 16'hfffe;
    LUT4 i1_4_lut_adj_43 (.A(n3047), .B(n28496), .C(n3048), .D(n3049), 
         .Z(n28578)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_43.init = 16'h8000;
    LUT4 i24570_2_lut_rep_184 (.A(n28522), .B(n13614), .Z(n38189)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24570_2_lut_rep_184.init = 16'heeee;
    LUT4 i24542_4_lut (.A(n3051), .B(n3050), .C(n28190), .D(n3052), 
         .Z(n28496)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24542_4_lut.init = 16'heccc;
    CCU2C add_26228_25 (.A0(n72_adj_5), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n69_adj_6), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30526), .COUT(n30527), .S0(n38[23]), .S1(n38[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_25.INIT0 = 16'h5550;
    defparam add_26228_25.INIT1 = 16'h5550;
    defparam add_26228_25.INJECT1_0 = "NO";
    defparam add_26228_25.INJECT1_1 = "NO";
    LUT4 i24238_3_lut (.A(n346), .B(n3053), .C(n3054), .Z(n28190)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24238_3_lut.init = 16'hecec;
    LUT4 div_13_i1866_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[14]), 
         .D(n2749), .Z(n2848_adj_646)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1866_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1869_3_lut_4_lut (.A(n28468), .B(n13622), .C(n2798[11]), 
         .D(n2752), .Z(n2851_adj_647)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1869_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_44 (.A(n2732_adj_648), .B(n2798_adj_2165[31]), 
         .C(n38239), .D(n2836), .Z(n35428)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_44.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_45 (.A(n2734_adj_650), .B(n2798_adj_2166[29]), 
         .C(n38240), .D(n2832), .Z(n36188)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_45.init = 16'hffca;
    PFUMX pwm_cnt_14__I_0_54_i24 (.BLUT(n16_adj_652), .ALUT(n22_adj_653), 
          .C0(n36752), .Z(n24_adj_654)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    LUT4 div_13_i2143_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[5]), 
         .D(n3154_adj_656), .Z(n3253_adj_657)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2143_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_26228_23 (.A0(n78_adj_7), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n75_adj_8), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30525), .COUT(n30526), .S0(n38[21]), .S1(n38[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_23.INIT0 = 16'h5550;
    defparam add_26228_23.INIT1 = 16'h5550;
    defparam add_26228_23.INJECT1_0 = "NO";
    defparam add_26228_23.INJECT1_1 = "NO";
    LUT4 div_13_i2127_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[21]), 
         .D(n3138_adj_661), .Z(n3237_adj_662)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_46 (.A(n2736_adj_663), .B(n2798_adj_2166[27]), 
         .C(n38240), .D(n2839_adj_665), .Z(n36196)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_46.init = 16'hffca;
    LUT4 div_13_i2144_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[4]), 
         .D(n347_adj_667), .Z(n3254_adj_668)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2144_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_47 (.A(n2646), .B(n2699[18]), .C(n38234), 
         .D(n2738), .Z(n35376)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_47.init = 16'hffca;
    CCU2C div_9_add_1445_5 (.A0(n13605), .B0(n28263), .C0(n2105[17]), 
          .D0(n2053), .A1(n13605), .B1(n28263), .C1(n2105[18]), .D1(n2052), 
          .CIN(n30672), .COUT(n30673), .S0(n2204[17]), .S1(n2204[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1445_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1445_5.INJECT1_0 = "NO";
    defparam div_9_add_1445_5.INJECT1_1 = "NO";
    LUT4 rem_10_mux_3_i9_3_lut_4_lut_4_lut (.A(n66_adj_9), .B(n38331), .C(n2[8]), 
         .D(n5), .Z(n592)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i9_3_lut_4_lut_4_lut.init = 16'hc088;
    LUT4 div_13_i2141_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[7]), 
         .D(n3152_adj_671), .Z(n3251_adj_672)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2141_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2126_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[22]), 
         .D(n3137_adj_674), .Z(n3236_adj_675)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1857_i7_3_lut_4_lut_4_lut (.A(n66_adj_9), .B(n38331), .C(n35[8]), 
         .D(n5), .Z(n343_adj_677)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i7_3_lut_4_lut_4_lut.init = 16'hc088;
    LUT4 i23479_2_lut_rep_317 (.A(n63_adj_10), .B(n3), .Z(n38322)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23479_2_lut_rep_317.init = 16'heeee;
    LUT4 div_13_i2120_3_lut_rep_177_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[28]), 
         .D(n3131), .Z(n38182)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2120_3_lut_rep_177_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1445_3 (.A0(n13605), .B0(n28263), .C0(n2105[15]), 
          .D0(n336), .A1(n13605), .B1(n28263), .C1(n2105[16]), .D1(n2054), 
          .CIN(n30671), .COUT(n30672), .S0(n2204[15]), .S1(n2204[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1445_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1445_3.INJECT1_0 = "NO";
    defparam div_9_add_1445_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_48 (.A(n2641), .B(n2699[23]), .C(n38234), 
         .D(n2735), .Z(n35384)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_48.init = 16'hffca;
    LUT4 i24510_2_lut_rep_229 (.A(n28462), .B(n13624), .Z(n38234)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24510_2_lut_rep_229.init = 16'heeee;
    CCU2C rem_10_add_1378_19 (.A0(n13604), .B0(n28333), .C0(n2006[31]), 
          .D0(n1940), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30589), .S0(n2105_adj_2168[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1378_19.INIT1 = 16'h0000;
    defparam rem_10_add_1378_19.INJECT1_0 = "NO";
    defparam rem_10_add_1378_19.INJECT1_1 = "NO";
    LUT4 i23442_2_lut_3_lut (.A(n63_adj_10), .B(n3), .C(n27382), .Z(duty0_14__N_426[7])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23442_2_lut_3_lut.init = 16'he0e0;
    LUT4 div_13_i2118_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[30]), 
         .D(n38192), .Z(n3228_adj_682)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1790_3_lut_rep_228_4_lut (.A(n28462), .B(n13624), .C(n2699[23]), 
         .D(n2641), .Z(n38233)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1790_3_lut_rep_228_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1797_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[16]), 
         .D(n2648), .Z(n2747)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2131_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[17]), 
         .D(n3142_adj_684), .Z(n3241_adj_685)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2131_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2124_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[24]), 
         .D(n3135_adj_687), .Z(n3234_adj_688)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1804_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[9]), 
         .D(n342), .Z(n2754)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1804_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1791_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[22]), 
         .D(n2642), .Z(n2741)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1791_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1713_19 (.A0(n13627), .B0(n28446), .C0(n2501[27]), 
          .D0(n2439), .A1(n13627), .B1(n28446), .C1(n2501[28]), .D1(n2438), 
          .CIN(n30958), .COUT(n30959), .S0(n2600[27]), .S1(n2600[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_19.INJECT1_0 = "NO";
    defparam div_13_add_1713_19.INJECT1_1 = "NO";
    CCU2C div_9_add_1445_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n48), .D1(n35[14]), 
          .COUT(n30671), .S1(n2204[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1445_1.INIT0 = 16'h0000;
    defparam div_9_add_1445_1.INIT1 = 16'habef;
    defparam div_9_add_1445_1.INJECT1_0 = "NO";
    defparam div_9_add_1445_1.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_11 (.A0(n13548), .B0(n28578), .C0(n3095[13]), 
          .D0(n3047), .A1(n13548), .B1(n28578), .C1(n3095[14]), .D1(n3046), 
          .CIN(n30790), .COUT(n30791), .S0(n3194[13]), .S1(n3194[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_11.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_11.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_11.INJECT1_0 = "NO";
    defparam div_9_add_2115_11.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_9 (.A0(n13548), .B0(n28578), .C0(n3095[11]), 
          .D0(n3049), .A1(n13548), .B1(n28578), .C1(n3095[12]), .D1(n3048), 
          .CIN(n30789), .COUT(n30790), .S0(n3194[11]), .S1(n3194[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_9.INIT0 = 16'hf1e0;
    defparam div_9_add_2115_9.INIT1 = 16'hf1e0;
    defparam div_9_add_2115_9.INJECT1_0 = "NO";
    defparam div_9_add_2115_9.INJECT1_1 = "NO";
    CCU2C div_9_add_2115_7 (.A0(n13548), .B0(n28578), .C0(n3095[9]), .D0(n3051), 
          .A1(n13548), .B1(n28578), .C1(n3095[10]), .D1(n3050), .CIN(n30788), 
          .COUT(n30789), .S0(n3194[9]), .S1(n3194[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_7.INIT0 = 16'h0e1f;
    defparam div_9_add_2115_7.INIT1 = 16'hf1e0;
    defparam div_9_add_2115_7.INJECT1_0 = "NO";
    defparam div_9_add_2115_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1713_17 (.A0(n13627), .B0(n28446), .C0(n2501[25]), 
          .D0(n2441), .A1(n13627), .B1(n28446), .C1(n2501[26]), .D1(n38255), 
          .CIN(n30957), .COUT(n30958), .S0(n2600[25]), .S1(n2600[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_17.INJECT1_0 = "NO";
    defparam div_13_add_1713_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_1177_15 (.A0(n38306), .B0(GND_net), .C0(n1709[30]), 
          .D0(GND_net), .A1(n38306), .B1(GND_net), .C1(n1709[31]), .D1(GND_net), 
          .CIN(n30669), .S0(n1808[30]), .S1(n1808[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1177_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1177_15.INJECT1_0 = "NO";
    defparam rem_10_add_1177_15.INJECT1_1 = "NO";
    LUT4 div_13_i1792_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[21]), 
         .D(n2643), .Z(n2742)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1792_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2115_5 (.A0(n13548), .B0(n28578), .C0(n3095[7]), .D0(n3053), 
          .A1(n13548), .B1(n28578), .C1(n3095[8]), .D1(n3052), .CIN(n30787), 
          .COUT(n30788), .S0(n3194[7]), .S1(n3194[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_5.INIT0 = 16'hf1e0;
    defparam div_9_add_2115_5.INIT1 = 16'hf1e0;
    defparam div_9_add_2115_5.INJECT1_0 = "NO";
    defparam div_9_add_2115_5.INJECT1_1 = "NO";
    LUT4 div_13_i2133_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[15]), 
         .D(n3144_adj_691), .Z(n3243_adj_692)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2133_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1796_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[17]), 
         .D(n2647), .Z(n2746)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1796_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1784_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[29]), 
         .D(n2635), .Z(n2734)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1784_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1794_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[19]), 
         .D(n2645), .Z(n2744)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1794_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2138_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[10]), 
         .D(n3149_adj_694), .Z(n3248_adj_695)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2138_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2115_3 (.A0(n13548), .B0(n28578), .C0(n3095[5]), .D0(n346), 
          .A1(n13548), .B1(n28578), .C1(n3095[6]), .D1(n3054), .CIN(n30786), 
          .COUT(n30787), .S0(n3194[5]), .S1(n3194[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_3.INIT0 = 16'hf1e0;
    defparam div_9_add_2115_3.INIT1 = 16'h0e1f;
    defparam div_9_add_2115_3.INJECT1_0 = "NO";
    defparam div_9_add_2115_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1713_15 (.A0(n13627), .B0(n28446), .C0(n2501[23]), 
          .D0(n2443), .A1(n13627), .B1(n28446), .C1(n2501[24]), .D1(n2442), 
          .CIN(n30956), .COUT(n30957), .S0(n2600[23]), .S1(n2600[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_15.INJECT1_0 = "NO";
    defparam div_13_add_1713_15.INJECT1_1 = "NO";
    LUT4 div_13_i2139_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[9]), 
         .D(n3150_adj_697), .Z(n3249_adj_698)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2139_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2115_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[4]), .D1(duty0_14__N_426[2]), 
          .COUT(n30786), .S1(n3194[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2115_1.INIT0 = 16'h0000;
    defparam div_9_add_2115_1.INIT1 = 16'h04bf;
    defparam div_9_add_2115_1.INJECT1_0 = "NO";
    defparam div_9_add_2115_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1713_13 (.A0(n13627), .B0(n28446), .C0(n2501[21]), 
          .D0(n2445), .A1(n13627), .B1(n28446), .C1(n2501[22]), .D1(n2444), 
          .CIN(n30955), .COUT(n30956), .S0(n2600[21]), .S1(n2600[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_13.INJECT1_0 = "NO";
    defparam div_13_add_1713_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_17 (.A0(n13604), .B0(n28333), .C0(n2006[29]), 
          .D0(n1942), .A1(n13604), .B1(n28333), .C1(n2006[30]), .D1(n1941), 
          .CIN(n30588), .COUT(n30589), .S0(n2105_adj_2168[29]), .S1(n2105_adj_2168[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1378_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1378_17.INJECT1_0 = "NO";
    defparam rem_10_add_1378_17.INJECT1_1 = "NO";
    CCU2C add_26228_21 (.A0(n84), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n81_adj_11), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n30524), .COUT(n30525), .S0(n38[19]), .S1(n38[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_21.INIT0 = 16'h5550;
    defparam add_26228_21.INIT1 = 16'h5550;
    defparam add_26228_21.INJECT1_0 = "NO";
    defparam add_26228_21.INJECT1_1 = "NO";
    CCU2C div_13_add_1713_11 (.A0(n13627), .B0(n28446), .C0(n2501[19]), 
          .D0(n2447), .A1(n13627), .B1(n28446), .C1(n2501[20]), .D1(n2446), 
          .CIN(n30954), .COUT(n30955), .S0(n2600[19]), .S1(n2600[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_11.INJECT1_0 = "NO";
    defparam div_13_add_1713_11.INJECT1_1 = "NO";
    LUT4 div_13_i2140_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[8]), 
         .D(n3151), .Z(n3250_adj_704)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2140_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1177_13 (.A0(n38306), .B0(GND_net), .C0(n1709[28]), 
          .D0(n38306), .A1(n38306), .B1(GND_net), .C1(n1709[29]), .D1(GND_net), 
          .CIN(n30668), .COUT(n30669), .S0(n1808[28]), .S1(n1808[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1177_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1177_13.INJECT1_0 = "NO";
    defparam rem_10_add_1177_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1713_9 (.A0(n13627), .B0(n28446), .C0(n2501[17]), 
          .D0(n2449), .A1(n13627), .B1(n28446), .C1(n2501[18]), .D1(n2448), 
          .CIN(n30953), .COUT(n30954), .S0(n2600[17]), .S1(n2600[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1713_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1713_9.INJECT1_0 = "NO";
    defparam div_13_add_1713_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1713_7 (.A0(n13627), .B0(n28446), .C0(n2501[15]), 
          .D0(n2451), .A1(n13627), .B1(n28446), .C1(n2501[16]), .D1(n2450), 
          .CIN(n30952), .COUT(n30953), .S0(n2600[15]), .S1(n2600[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1713_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1713_7.INJECT1_0 = "NO";
    defparam div_13_add_1713_7.INJECT1_1 = "NO";
    LUT4 div_13_i1782_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[31]), 
         .D(n38241), .Z(n2732)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1782_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1798_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[15]), 
         .D(n2649), .Z(n2748)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1798_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2048_27 (.A0(n13549), .B0(n28574), .C0(n2996[30]), 
          .D0(n2931), .A1(n13549), .B1(n28574), .C1(n2996[31]), .D1(n2930_adj_706), 
          .CIN(n30784), .S0(n3095[30]), .S1(n3095[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_27.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_27.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_27.INJECT1_0 = "NO";
    defparam div_9_add_2048_27.INJECT1_1 = "NO";
    LUT4 div_13_i1795_3_lut_rep_227_4_lut (.A(n28462), .B(n13624), .C(n2699[18]), 
         .D(n2646), .Z(n38232)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1795_3_lut_rep_227_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1177_11 (.A0(n38306), .B0(GND_net), .C0(n1709[26]), 
          .D0(GND_net), .A1(n38306), .B1(GND_net), .C1(n1709[27]), .D1(GND_net), 
          .CIN(n30667), .COUT(n30668), .S0(n1808[26]), .S1(n1808[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_11.INIT0 = 16'hf1e0;
    defparam rem_10_add_1177_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1177_11.INJECT1_0 = "NO";
    defparam rem_10_add_1177_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_15 (.A0(n13604), .B0(n28333), .C0(n2006[27]), 
          .D0(n1944), .A1(n13604), .B1(n28333), .C1(n2006[28]), .D1(n1943), 
          .CIN(n30587), .COUT(n30588), .S0(n2105_adj_2168[27]), .S1(n2105_adj_2168[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1378_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1378_15.INJECT1_0 = "NO";
    defparam rem_10_add_1378_15.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_25 (.A0(n13549), .B0(n28574), .C0(n2996[28]), 
          .D0(n38221), .A1(n13549), .B1(n28574), .C1(n2996[29]), .D1(n2932_adj_709), 
          .CIN(n30783), .COUT(n30784), .S0(n3095[28]), .S1(n3095[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_25.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_25.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_25.INJECT1_0 = "NO";
    defparam div_9_add_2048_25.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_23 (.A0(n13549), .B0(n28574), .C0(n2996[26]), 
          .D0(n2935_adj_710), .A1(n13549), .B1(n28574), .C1(n2996[27]), 
          .D1(n2934_adj_711), .CIN(n30782), .COUT(n30783), .S0(n3095[26]), 
          .S1(n3095[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_23.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_23.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_23.INJECT1_0 = "NO";
    defparam div_9_add_2048_23.INJECT1_1 = "NO";
    CCU2C rem_10_add_1177_9 (.A0(n38306), .B0(GND_net), .C0(n1709[24]), 
          .D0(GND_net), .A1(n38306), .B1(GND_net), .C1(n1709[25]), .D1(n38306), 
          .CIN(n30666), .COUT(n30667), .S0(n1808[24]), .S1(n1808[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1177_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1177_9.INJECT1_0 = "NO";
    defparam rem_10_add_1177_9.INJECT1_1 = "NO";
    LUT4 div_13_i1787_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[26]), 
         .D(n2638), .Z(n2737)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1787_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2410_3_lut_4_lut (.A(n28462), .B(n13624), .C(n3556), 
         .D(n4990[8]), .Z(n197[8])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2410_3_lut_4_lut.init = 16'hfe0e;
    CCU2C div_13_add_1713_5 (.A0(n13627), .B0(n28446), .C0(n2501[13]), 
          .D0(n2453), .A1(n13627), .B1(n28446), .C1(n2501[14]), .D1(n2452), 
          .CIN(n30951), .COUT(n30952), .S0(n2600[13]), .S1(n2600[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1713_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1713_5.INJECT1_0 = "NO";
    defparam div_13_add_1713_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_13 (.A0(n13604), .B0(n28333), .C0(n2006[25]), 
          .D0(n1946), .A1(n13604), .B1(n28333), .C1(n2006[26]), .D1(n1945), 
          .CIN(n30586), .COUT(n30587), .S0(n2105_adj_2168[25]), .S1(n2105_adj_2168[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1378_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1378_13.INJECT1_0 = "NO";
    defparam rem_10_add_1378_13.INJECT1_1 = "NO";
    CCU2C add_26228_19 (.A0(n90), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n87), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30523), 
          .COUT(n30524), .S0(n38[17]), .S1(n38[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_19.INIT0 = 16'h5550;
    defparam add_26228_19.INIT1 = 16'h5550;
    defparam add_26228_19.INJECT1_0 = "NO";
    defparam add_26228_19.INJECT1_1 = "NO";
    LUT4 div_13_i2142_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[6]), 
         .D(n3153_adj_717), .Z(n3252_adj_718)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2142_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2202_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[13]), 
         .D(n3245_adj_720), .Z(n3344_adj_721)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2202_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2119_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[29]), 
         .D(n38193), .Z(n3229_adj_723)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1123_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[20]), 
         .D(n331), .Z(n1753_adj_724)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1785_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[28]), 
         .D(n2636), .Z(n2735)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1785_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1713_3 (.A0(n13627), .B0(n28446), .C0(n2501[11]), 
          .D0(n340), .A1(n13627), .B1(n28446), .C1(n2501[12]), .D1(n2454), 
          .CIN(n30950), .COUT(n30951), .S0(n2600[11]), .S1(n2600[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1713_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1713_3.INJECT1_0 = "NO";
    defparam div_13_add_1713_3.INJECT1_1 = "NO";
    LUT4 div_13_i1800_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[13]), 
         .D(n2651), .Z(n2750)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1800_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2117_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[31]), 
         .D(n3128), .Z(n3227_adj_726)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2117_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1713_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n341_adj_605), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30950), .S1(n2600[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1713_1.INIT0 = 16'h0000;
    defparam div_13_add_1713_1.INIT1 = 16'h555a;
    defparam div_13_add_1713_1.INJECT1_0 = "NO";
    defparam div_13_add_1713_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_11 (.A0(n13604), .B0(n28333), .C0(n2006[23]), 
          .D0(n1948), .A1(n13604), .B1(n28333), .C1(n2006[24]), .D1(n1947), 
          .CIN(n30585), .COUT(n30586), .S0(n2105_adj_2168[23]), .S1(n2105_adj_2168[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_11.INIT0 = 16'hf1e0;
    defparam rem_10_add_1378_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1378_11.INJECT1_0 = "NO";
    defparam rem_10_add_1378_11.INJECT1_1 = "NO";
    LUT4 div_13_i2130_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[18]), 
         .D(n3141_adj_730), .Z(n3240_adj_564)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2130_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1799_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[14]), 
         .D(n2650), .Z(n2749)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1799_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1646_21 (.A0(n13630), .B0(n28442), .C0(n2402[30]), 
          .D0(n2337), .A1(n13630), .B1(n28442), .C1(n2402[31]), .D1(n2336), 
          .CIN(n30948), .S0(n2501[30]), .S1(n2501[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_21.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_21.INJECT1_0 = "NO";
    defparam div_13_add_1646_21.INJECT1_1 = "NO";
    CCU2C rem_10_add_1177_7 (.A0(n38306), .B0(GND_net), .C0(n1709[22]), 
          .D0(n38306), .A1(n38306), .B1(GND_net), .C1(n1709[23]), .D1(GND_net), 
          .CIN(n30665), .COUT(n30666), .S0(n1808[22]), .S1(n1808[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_7.INIT0 = 16'hf1e0;
    defparam rem_10_add_1177_7.INIT1 = 16'h0e1f;
    defparam rem_10_add_1177_7.INJECT1_0 = "NO";
    defparam rem_10_add_1177_7.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_9 (.A0(n13604), .B0(n28333), .C0(n2006[21]), 
          .D0(n1950), .A1(n13604), .B1(n28333), .C1(n2006[22]), .D1(n1949), 
          .CIN(n30584), .COUT(n30585), .S0(n2105_adj_2168[21]), .S1(n2105_adj_2168[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1378_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1378_9.INJECT1_0 = "NO";
    defparam rem_10_add_1378_9.INJECT1_1 = "NO";
    LUT4 div_13_i2132_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[16]), 
         .D(n3143), .Z(n3242_adj_603)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2132_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1788_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[25]), 
         .D(n2639), .Z(n2738)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1788_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1177_5 (.A0(n38306), .B0(GND_net), .C0(n1709[20]), 
          .D0(n38306), .A1(n38306), .B1(GND_net), .C1(n1709[21]), .D1(n38306), 
          .CIN(n30664), .COUT(n30665), .S0(n1808[20]), .S1(n1808[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_5.INIT0 = 16'h0e1f;
    defparam rem_10_add_1177_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1177_5.INJECT1_0 = "NO";
    defparam rem_10_add_1177_5.INJECT1_1 = "NO";
    LUT4 div_13_i2203_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[12]), 
         .D(n3246_adj_736), .Z(n3345_adj_634)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2203_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1802_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[11]), 
         .D(n2653), .Z(n2752)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1802_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32161_4_lut (.A(n38392), .B(n38391), .C(n38390), .D(n36852), 
         .Z(n36866)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32161_4_lut.init = 16'hfffe;
    LUT4 div_13_i1783_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[30]), 
         .D(n2634), .Z(n2733)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1783_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_2048_21 (.A0(n13549), .B0(n28574), .C0(n2996[24]), 
          .D0(n2937), .A1(n13549), .B1(n28574), .C1(n2996[25]), .D1(n2936_adj_737), 
          .CIN(n30781), .COUT(n30782), .S0(n3095[24]), .S1(n3095[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_21.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_21.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_21.INJECT1_0 = "NO";
    defparam div_9_add_2048_21.INJECT1_1 = "NO";
    LUT4 div_13_i1789_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[24]), 
         .D(n2640), .Z(n2739)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1789_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1378_7 (.A0(n13604), .B0(n28333), .C0(n2006[19]), 
          .D0(n1952), .A1(n13604), .B1(n28333), .C1(n2006[20]), .D1(n1951), 
          .CIN(n30583), .COUT(n30584), .S0(n2105_adj_2168[19]), .S1(n2105_adj_2168[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_7.INIT0 = 16'hf1e0;
    defparam rem_10_add_1378_7.INIT1 = 16'h0e1f;
    defparam rem_10_add_1378_7.INJECT1_0 = "NO";
    defparam rem_10_add_1378_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1646_19 (.A0(n13630), .B0(n28442), .C0(n2402[28]), 
          .D0(n2339), .A1(n13630), .B1(n28442), .C1(n2402[29]), .D1(n2338), 
          .CIN(n30947), .COUT(n30948), .S0(n2501[28]), .S1(n2501[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_19.INJECT1_0 = "NO";
    defparam div_13_add_1646_19.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_49 (.A(n35556), .B(n2444), .C(n35540), .D(n2445), 
         .Z(n13627)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_49.init = 16'hfffe;
    CCU2C div_9_add_2048_19 (.A0(n13549), .B0(n28574), .C0(n2996[22]), 
          .D0(n2939_adj_740), .A1(n13549), .B1(n28574), .C1(n2996[23]), 
          .D1(n2938_adj_741), .CIN(n30780), .COUT(n30781), .S0(n3095[22]), 
          .S1(n3095[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_19.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_19.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_19.INJECT1_0 = "NO";
    defparam div_9_add_2048_19.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_17 (.A0(n13549), .B0(n28574), .C0(n2996[20]), 
          .D0(n2941), .A1(n13549), .B1(n28574), .C1(n2996[21]), .D1(n2940_adj_742), 
          .CIN(n30779), .COUT(n30780), .S0(n3095[20]), .S1(n3095[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_17.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_17.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_17.INJECT1_0 = "NO";
    defparam div_9_add_2048_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_50 (.A(n2438), .B(n35552), .C(n35538), .D(n2441), 
         .Z(n35556)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_50.init = 16'hfffe;
    CCU2C rem_10_add_1378_5 (.A0(n13604), .B0(n28333), .C0(n2006[17]), 
          .D0(n1954), .A1(n13604), .B1(n28333), .C1(n2006[18]), .D1(n1953), 
          .CIN(n30582), .COUT(n30583), .S0(n2105_adj_2168[17]), .S1(n2105_adj_2168[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_5.INIT0 = 16'h0e1f;
    defparam rem_10_add_1378_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1378_5.INJECT1_0 = "NO";
    defparam rem_10_add_1378_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_51 (.A(n2443), .B(n2437), .C(n2446), .D(n2439), 
         .Z(n35552)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_51.init = 16'hfffe;
    LUT4 div_13_i1803_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[10]), 
         .D(n2654), .Z(n2753)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1803_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_52 (.A(n2448), .B(n28309), .C(n2447), .D(n2449), 
         .Z(n28446)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_52.init = 16'h8000;
    LUT4 i24356_4_lut (.A(n2451), .B(n2450), .C(n28052), .D(n2452), 
         .Z(n28309)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24356_4_lut.init = 16'heccc;
    CCU2C div_9_add_2048_15 (.A0(n13549), .B0(n28574), .C0(n2996[18]), 
          .D0(n2943_adj_745), .A1(n13549), .B1(n28574), .C1(n2996[19]), 
          .D1(n2942_adj_746), .CIN(n30778), .COUT(n30779), .S0(n3095[18]), 
          .S1(n3095[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_15.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_15.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_15.INJECT1_0 = "NO";
    defparam div_9_add_2048_15.INJECT1_1 = "NO";
    LUT4 div_13_i1793_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[20]), 
         .D(n2644), .Z(n2743)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1793_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1646_17 (.A0(n13630), .B0(n28442), .C0(n2402[26]), 
          .D0(n2341), .A1(n13630), .B1(n28442), .C1(n2402[27]), .D1(n2340), 
          .CIN(n30946), .COUT(n30947), .S0(n2501[26]), .S1(n2501[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_17.INJECT1_0 = "NO";
    defparam div_13_add_1646_17.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_13 (.A0(n13549), .B0(n28574), .C0(n2996[16]), 
          .D0(n2945_adj_747), .A1(n13549), .B1(n28574), .C1(n2996[17]), 
          .D1(n2944_adj_748), .CIN(n30777), .COUT(n30778), .S0(n3095[16]), 
          .S1(n3095[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_13.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_13.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_13.INJECT1_0 = "NO";
    defparam div_9_add_2048_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1177_3 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[18]), 
          .A1(n38307), .B1(n1709[19]), .C1(n2[19]), .D1(n38306), .CIN(n30663), 
          .COUT(n30664), .S0(n1808[18]), .S1(n1808[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_3.INIT0 = 16'h2000;
    defparam rem_10_add_1177_3.INIT1 = 16'hcca0;
    defparam rem_10_add_1177_3.INJECT1_0 = "NO";
    defparam rem_10_add_1177_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1646_15 (.A0(n13630), .B0(n28442), .C0(n2402[24]), 
          .D0(n38262), .A1(n13630), .B1(n28442), .C1(n2402[25]), .D1(n2342), 
          .CIN(n30945), .COUT(n30946), .S0(n2501[24]), .S1(n2501[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_15.INJECT1_0 = "NO";
    defparam div_13_add_1646_15.INJECT1_1 = "NO";
    CCU2C add_26228_17 (.A0(n96), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n93), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30522), 
          .COUT(n30523), .S0(n38[15]), .S1(n38[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_17.INIT0 = 16'h5550;
    defparam add_26228_17.INIT1 = 16'h5550;
    defparam add_26228_17.INJECT1_0 = "NO";
    defparam add_26228_17.INJECT1_1 = "NO";
    LUT4 div_13_i2121_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[27]), 
         .D(n38194), .Z(n3231_adj_612)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24102_3_lut (.A(n340), .B(n2453), .C(n2454), .Z(n28052)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24102_3_lut.init = 16'hecec;
    CCU2C rem_10_add_1177_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n39), .D1(n2[17]), 
          .COUT(n30663));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1177_1.INIT0 = 16'h000F;
    defparam rem_10_add_1177_1.INIT1 = 16'habef;
    defparam rem_10_add_1177_1.INJECT1_0 = "NO";
    defparam rem_10_add_1177_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1646_13 (.A0(n13630), .B0(n28442), .C0(n2402[22]), 
          .D0(n2345), .A1(n13630), .B1(n28442), .C1(n2402[23]), .D1(n2344), 
          .CIN(n30944), .COUT(n30945), .S0(n2501[22]), .S1(n2501[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_13.INJECT1_0 = "NO";
    defparam div_13_add_1646_13.INJECT1_1 = "NO";
    LUT4 div_13_i1786_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[27]), 
         .D(n2637), .Z(n2736)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1786_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2128_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[20]), 
         .D(n3139_adj_753), .Z(n3238_adj_754)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2128_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1378_17 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[30]), 
          .D0(n1941_adj_756), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[31]), 
          .D1(n1940_adj_758), .CIN(n30661), .S0(n2105[30]), .S1(n2105[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1378_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1378_17.INJECT1_0 = "NO";
    defparam div_9_add_1378_17.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_11 (.A0(n13549), .B0(n28574), .C0(n2996[14]), 
          .D0(n2947), .A1(n13549), .B1(n28574), .C1(n2996[15]), .D1(n2946_adj_759), 
          .CIN(n30776), .COUT(n30777), .S0(n3095[14]), .S1(n3095[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_11.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_11.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_11.INJECT1_0 = "NO";
    defparam div_9_add_2048_11.INJECT1_1 = "NO";
    LUT4 div_13_i1801_3_lut_4_lut (.A(n28462), .B(n13624), .C(n2699[12]), 
         .D(n2652), .Z(n2751)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1801_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_53 (.A(n2738_adj_760), .B(n2798_adj_2165[25]), 
         .C(n38239), .D(n2839), .Z(n35424)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_53.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_54 (.A(n2742_adj_762), .B(n2798_adj_2166[21]), 
         .C(n38240), .D(n2842_adj_764), .Z(n36186)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_54.init = 16'hffca;
    LUT4 div_13_i2416_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3556), 
         .D(n4990[2]), .Z(n197[2])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2416_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i24596_2_lut_rep_172 (.A(n28512), .B(n13602), .Z(n38177)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24596_2_lut_rep_172.init = 16'heeee;
    LUT4 div_13_i2122_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[26]), 
         .D(n3133), .Z(n3232_adj_766)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2135_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[13]), 
         .D(n3146_adj_768), .Z(n3245_adj_720)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2135_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2136_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[12]), 
         .D(n3147_adj_770), .Z(n3246_adj_736)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2136_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2129_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[19]), 
         .D(n3140_adj_772), .Z(n3239_adj_773)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2129_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_55 (.A(n2753_adj_774), .B(n2798_adj_2165[10]), 
         .C(n38239), .D(n2851), .Z(n34684)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_55.init = 16'hca00;
    CCU2C div_13_add_1646_11 (.A0(n13630), .B0(n28442), .C0(n2402[20]), 
          .D0(n2347), .A1(n13630), .B1(n28442), .C1(n2402[21]), .D1(n2346), 
          .CIN(n30943), .COUT(n30944), .S0(n2501[20]), .S1(n2501[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_11.INJECT1_0 = "NO";
    defparam div_13_add_1646_11.INJECT1_1 = "NO";
    LUT4 div_13_i2415_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3556), 
         .D(n4990[3]), .Z(n197[3])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2415_3_lut_4_lut.init = 16'hfe0e;
    CCU2C div_9_add_1378_15 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[28]), 
          .D0(n1943_adj_777), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[29]), 
          .D1(n1942_adj_779), .CIN(n30660), .COUT(n30661), .S0(n2105[28]), 
          .S1(n2105[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1378_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1378_15.INJECT1_0 = "NO";
    defparam div_9_add_1378_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_56 (.A(n2741_adj_780), .B(n2798_adj_2165[22]), 
         .C(n38239), .D(n2844), .Z(n35434)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_56.init = 16'hffca;
    CCU2C div_9_add_1378_13 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[26]), 
          .D0(n1945_adj_783), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[27]), 
          .D1(n1944_adj_785), .CIN(n30659), .COUT(n30660), .S0(n2105[26]), 
          .S1(n2105[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1378_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1378_13.INJECT1_0 = "NO";
    defparam div_9_add_1378_13.INJECT1_1 = "NO";
    LUT4 n3395_bdd_4_lut_32316 (.A(n3392[29]), .B(n3392[24]), .C(n3392[19]), 
         .D(n3392[13]), .Z(n37667)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3395_bdd_4_lut_32316.init = 16'hfffe;
    LUT4 i24500_2_lut_rep_234 (.A(n28373), .B(n13626), .Z(n38239)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24500_2_lut_rep_234.init = 16'heeee;
    LUT4 i32183_4_lut (.A(n38386), .B(n38385), .C(n38384), .D(n36795), 
         .Z(n36809)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i32183_4_lut.init = 16'hfffe;
    CCU2C div_9_add_2048_9 (.A0(n13549), .B0(n28574), .C0(n2996[12]), 
          .D0(n2949_adj_786), .A1(n13549), .B1(n28574), .C1(n2996[13]), 
          .D1(n2948_adj_787), .CIN(n30775), .COUT(n30776), .S0(n3095[12]), 
          .S1(n3095[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_9.INIT0 = 16'hf1e0;
    defparam div_9_add_2048_9.INIT1 = 16'hf1e0;
    defparam div_9_add_2048_9.INJECT1_0 = "NO";
    defparam div_9_add_2048_9.INJECT1_1 = "NO";
    CCU2C add_26228_15 (.A0(n102), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n99), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30521), 
          .COUT(n30522), .S0(n38[13]), .S1(n38[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_15.INIT0 = 16'h5550;
    defparam add_26228_15.INIT1 = 16'h5550;
    defparam add_26228_15.INJECT1_0 = "NO";
    defparam add_26228_15.INJECT1_1 = "NO";
    LUT4 rem_10_i1849_3_lut_rep_224_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[31]), 
         .D(n2732_adj_648), .Z(n38229)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1849_3_lut_rep_224_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1855_3_lut_rep_230_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[25]), 
         .D(n2738_adj_760), .Z(n38235)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1855_3_lut_rep_230_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1870_3_lut_rep_232_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[10]), 
         .D(n2753_adj_774), .Z(n38237)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1870_3_lut_rep_232_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1858_3_lut_rep_233_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[22]), 
         .D(n2741_adj_780), .Z(n38238)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1858_3_lut_rep_233_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_57 (.A(n27382), .B(n3), .C(n54), .Z(duty0_14__N_426[10])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_57.init = 16'h2020;
    LUT4 div_13_i2125_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[23]), 
         .D(n3136_adj_791), .Z(n3235_adj_792)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2123_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[25]), 
         .D(n3134_adj_794), .Z(n3233_adj_795)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1862_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[18]), 
         .D(n2745), .Z(n2844)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1862_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_326 (.A(n3), .B(n27382), .Z(n38331)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_326.init = 16'h4444;
    LUT4 rem_10_i1854_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[26]), 
         .D(n2737_adj_798), .Z(n2836)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1854_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1378_11 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[24]), 
          .D0(n1947_adj_800), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[25]), 
          .D1(n1946_adj_802), .CIN(n30658), .COUT(n30659), .S0(n2105[24]), 
          .S1(n2105[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1378_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1378_11.INJECT1_0 = "NO";
    defparam div_9_add_1378_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_3 (.A0(n12154), .B0(n5), .C0(n45), .D0(n2[15]), 
          .A1(n13604), .B1(n28333), .C1(n2006[16]), .D1(n584), .CIN(n30581), 
          .COUT(n30582), .S0(n2105_adj_2168[15]), .S1(n2105_adj_2168[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_3.INIT0 = 16'h5410;
    defparam rem_10_add_1378_3.INIT1 = 16'hf1e0;
    defparam rem_10_add_1378_3.INJECT1_0 = "NO";
    defparam rem_10_add_1378_3.INJECT1_1 = "NO";
    LUT4 div_13_i2134_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[14]), 
         .D(n3145_adj_806), .Z(n3244_adj_807)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2134_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2261_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[21]), 
         .D(n3336_adj_808), .Z(n43)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2261_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1646_9 (.A0(n13630), .B0(n28442), .C0(n2402[18]), 
          .D0(n2349), .A1(n13630), .B1(n28442), .C1(n2402[19]), .D1(n2348), 
          .CIN(n30942), .COUT(n30943), .S0(n2501[18]), .S1(n2501[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1646_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1646_9.INJECT1_0 = "NO";
    defparam div_13_add_1646_9.INJECT1_1 = "NO";
    LUT4 div_13_i2137_3_lut_4_lut (.A(n28522), .B(n13614), .C(n3194_adj_2167[11]), 
         .D(n3148_adj_810), .Z(n3247_adj_811)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2137_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1646_7 (.A0(n13630), .B0(n28442), .C0(n2402[16]), 
          .D0(n2351), .A1(n13630), .B1(n28442), .C1(n2402[17]), .D1(n2350), 
          .CIN(n30941), .COUT(n30942), .S0(n2501[16]), .S1(n2501[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1646_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1646_7.INJECT1_0 = "NO";
    defparam div_13_add_1646_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1646_5 (.A0(n13630), .B0(n28442), .C0(n2402[14]), 
          .D0(n2353), .A1(n13630), .B1(n28442), .C1(n2402[15]), .D1(n2352), 
          .CIN(n30940), .COUT(n30941), .S0(n2501[14]), .S1(n2501[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1646_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1646_5.INJECT1_0 = "NO";
    defparam div_13_add_1646_5.INJECT1_1 = "NO";
    CCU2C div_13_add_1646_3 (.A0(n13630), .B0(n28442), .C0(n2402[12]), 
          .D0(n339), .A1(n13630), .B1(n28442), .C1(n2402[13]), .D1(n2354), 
          .CIN(n30939), .COUT(n30940), .S0(n2501[12]), .S1(n2501[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1646_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1646_3.INJECT1_0 = "NO";
    defparam div_13_add_1646_3.INJECT1_1 = "NO";
    LUT4 div_9_i2255_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[27]), 
         .D(n3330_adj_812), .Z(n55)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2255_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32211_4_lut (.A(n38380), .B(n38379), .C(n38378), .D(n36738), 
         .Z(n36752)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i32211_4_lut.init = 16'hfffe;
    LUT4 rem_10_i1852_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[28]), 
         .D(n2735_adj_814), .Z(n2834)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1852_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1856_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[24]), 
         .D(n2739_adj_816), .Z(n2838_adj_525)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1856_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_58 (.A(n35742), .B(n1944), .C(n1941), .D(n1945), 
         .Z(n13604)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_58.init = 16'hfffe;
    LUT4 rem_10_i1863_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[17]), 
         .D(n2746_adj_818), .Z(n2845)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1863_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_59 (.A(n1942), .B(n1943), .C(n1940), .D(n1946), 
         .Z(n35742)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_59.init = 16'hfffe;
    LUT4 i1_4_lut_adj_60 (.A(n1947), .B(n28174), .C(n1948), .D(n1949), 
         .Z(n28333)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_60.init = 16'h8000;
    LUT4 i24222_4_lut (.A(n1951), .B(n1950), .C(n27898), .D(n1952), 
         .Z(n28174)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24222_4_lut.init = 16'heccc;
    LUT4 i23949_3_lut (.A(n584), .B(n1953), .C(n1954), .Z(n27898)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23949_3_lut.init = 16'hecec;
    LUT4 i23008_2_lut_rep_302_3_lut (.A(n3), .B(n27382), .C(n5), .Z(n38307)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i23008_2_lut_rep_302_3_lut.init = 16'h4040;
    CCU2C div_9_add_2048_7 (.A0(n13549), .B0(n28574), .C0(n2996[10]), 
          .D0(n2951_adj_819), .A1(n13549), .B1(n28574), .C1(n2996[11]), 
          .D1(n2950_adj_820), .CIN(n30774), .COUT(n30775), .S0(n3095[10]), 
          .S1(n3095[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_7.INIT0 = 16'h0e1f;
    defparam div_9_add_2048_7.INIT1 = 16'hf1e0;
    defparam div_9_add_2048_7.INJECT1_0 = "NO";
    defparam div_9_add_2048_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_61 (.A(n36154), .B(n36144), .C(n2943_adj_745), .D(n2938_adj_741), 
         .Z(n13549)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_61.init = 16'hfffe;
    LUT4 i1_4_lut_adj_62 (.A(n36148), .B(n36134), .C(n36146), .D(n2941), 
         .Z(n36154)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_62.init = 16'hfffe;
    LUT4 rem_10_i1861_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[19]), 
         .D(n2744_adj_822), .Z(n2843)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1861_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_63 (.A(n3130), .B(n3194[29]), .C(n38197), 
         .D(n3234), .Z(n36090)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_63.init = 16'hffca;
    LUT4 rem_10_i1864_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[16]), 
         .D(n2747_adj_824), .Z(n2846)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1864_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_64 (.A(n27382), .B(n3), .C(n51), .Z(duty0_14__N_426[11])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_64.init = 16'h2020;
    LUT4 rem_10_i1851_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[29]), 
         .D(n38242), .Z(n2833)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1851_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_65 (.A(n2944_adj_748), .B(n2934_adj_711), .C(n2946_adj_759), 
         .D(n2936_adj_737), .Z(n36144)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_65.init = 16'hfffe;
    LUT4 i1_4_lut_adj_66 (.A(n2935_adj_710), .B(n2937), .C(n2931), .D(n2932_adj_709), 
         .Z(n36148)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_66.init = 16'hfffe;
    CCU2C div_9_add_1378_9 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[22]), 
          .D0(n1949_adj_827), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[23]), 
          .D1(n1948_adj_829), .CIN(n30657), .COUT(n30658), .S0(n2105[22]), 
          .S1(n2105[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1378_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1378_9.INJECT1_0 = "NO";
    defparam div_9_add_1378_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_67 (.A(n2930_adj_706), .B(n2939_adj_740), .C(n2945_adj_747), 
         .D(n2940_adj_742), .Z(n36146)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_67.init = 16'hfffe;
    CCU2C div_9_add_2048_5 (.A0(n13549), .B0(n28574), .C0(n2996[8]), .D0(n2953_adj_830), 
          .A1(n13549), .B1(n28574), .C1(n2996[9]), .D1(n2952), .CIN(n30773), 
          .COUT(n30774), .S0(n3095[8]), .S1(n3095[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_5.INIT0 = 16'hf1e0;
    defparam div_9_add_2048_5.INIT1 = 16'hf1e0;
    defparam div_9_add_2048_5.INJECT1_0 = "NO";
    defparam div_9_add_2048_5.INJECT1_1 = "NO";
    LUT4 i9910_2_lut_3_lut_4_lut (.A(n3), .B(n27382), .C(n35[18]), .D(n5), 
         .Z(n333)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i9910_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_68 (.A(n2947), .B(n28502), .C(n2948_adj_787), .D(n2949_adj_786), 
         .Z(n28574)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_68.init = 16'h8000;
    LUT4 i24548_4_lut (.A(n2951_adj_819), .B(n2950_adj_820), .C(n28202), 
         .D(n2952), .Z(n28502)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24548_4_lut.init = 16'heccc;
    CCU2C div_9_add_1378_7 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[20]), 
          .D0(n1951_adj_833), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[21]), 
          .D1(n1950_adj_835), .CIN(n30656), .COUT(n30657), .S0(n2105[20]), 
          .S1(n2105[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1378_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1378_7.INJECT1_0 = "NO";
    defparam div_9_add_1378_7.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_3 (.A0(n13549), .B0(n28574), .C0(n2996[6]), .D0(n345), 
          .A1(n13549), .B1(n28574), .C1(n2996[7]), .D1(n2954_adj_836), 
          .CIN(n30772), .COUT(n30773), .S0(n3095[6]), .S1(n3095[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_3.INIT0 = 16'hf1e0;
    defparam div_9_add_2048_3.INIT1 = 16'h0e1f;
    defparam div_9_add_2048_3.INJECT1_0 = "NO";
    defparam div_9_add_2048_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1378_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n48), .D1(n2[14]), 
          .COUT(n30581));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1378_1.INIT0 = 16'h000F;
    defparam rem_10_add_1378_1.INIT1 = 16'habef;
    defparam rem_10_add_1378_1.INJECT1_0 = "NO";
    defparam rem_10_add_1378_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1378_5 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[18]), 
          .D0(n1953_adj_838), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[19]), 
          .D1(n1952_adj_840), .CIN(n30655), .COUT(n30656), .S0(n2105[18]), 
          .S1(n2105[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1378_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1378_5.INJECT1_0 = "NO";
    defparam div_9_add_1378_5.INJECT1_1 = "NO";
    LUT4 i24250_3_lut (.A(n345), .B(n2953_adj_830), .C(n2954_adj_836), 
         .Z(n28202)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24250_3_lut.init = 16'hecec;
    CCU2C div_13_add_1646_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n340), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30939), .S1(n2501[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1646_1.INIT0 = 16'h0000;
    defparam div_13_add_1646_1.INIT1 = 16'h555a;
    defparam div_13_add_1646_1.INJECT1_0 = "NO";
    defparam div_13_add_1646_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_69 (.A(n35624), .B(n2338), .C(n2337), .D(n2339), 
         .Z(n13630)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_69.init = 16'hfffe;
    PFUMX pwm_cnt_14__I_0_51_i28 (.BLUT(n12_adj_841), .ALUT(n26_adj_842), 
          .C0(n36947), .Z(n28)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    CCU2C div_13_add_1579_21 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[31]), 
          .D0(n2237), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30938), .S0(n2402[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_21.INIT1 = 16'h0000;
    defparam div_13_add_1579_21.INJECT1_0 = "NO";
    defparam div_13_add_1579_21.INJECT1_1 = "NO";
    LUT4 i9931_2_lut_rep_301_3_lut_4_lut (.A(n3), .B(n27382), .C(n2[19]), 
         .D(n5), .Z(n38306)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i9931_2_lut_rep_301_3_lut_4_lut.init = 16'h4000;
    LUT4 i9909_2_lut_rep_300_3_lut_4_lut (.A(n3), .B(n27382), .C(n35[19]), 
         .D(n5), .Z(n38305)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i9909_2_lut_rep_300_3_lut_4_lut.init = 16'h4000;
    LUT4 i23619_2_lut_rep_316_3_lut (.A(n3), .B(n27382), .C(n66_adj_9), 
         .Z(n38321)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i23619_2_lut_rep_316_3_lut.init = 16'h4040;
    CCU2C rem_10_add_1445_19 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[30]), 
          .D0(n2040_adj_844), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[31]), 
          .D1(n2039_adj_845), .CIN(n30579), .S0(n2204_adj_2172[30]), .S1(n2204_adj_2172[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1445_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1445_19.INJECT1_0 = "NO";
    defparam rem_10_add_1445_19.INJECT1_1 = "NO";
    CCU2C div_9_add_2048_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n75_adj_1), .D1(n35[5]), 
          .COUT(n30772), .S1(n3095[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2048_1.INIT0 = 16'h0000;
    defparam div_9_add_2048_1.INIT1 = 16'habef;
    defparam div_9_add_2048_1.INJECT1_0 = "NO";
    defparam div_9_add_2048_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1445_17 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[28]), 
          .D0(n2042_adj_849), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[29]), 
          .D1(n2041_adj_850), .CIN(n30578), .COUT(n30579), .S0(n2204_adj_2172[28]), 
          .S1(n2204_adj_2172[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1445_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1445_17.INJECT1_0 = "NO";
    defparam rem_10_add_1445_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_70 (.A(n2346), .B(n35620), .C(n35608), .D(n2340), 
         .Z(n35624)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_70.init = 16'hfffe;
    LUT4 i23486_2_lut_rep_327 (.A(n69_adj_12), .B(n3), .Z(n38332)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23486_2_lut_rep_327.init = 16'heeee;
    CCU2C div_13_add_1579_19 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[29]), 
          .D0(n2239), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[30]), 
          .D1(n2238), .CIN(n30937), .COUT(n30938), .S0(n2402[29]), .S1(n2402[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1579_19.INJECT1_0 = "NO";
    defparam div_13_add_1579_19.INJECT1_1 = "NO";
    CCU2C div_9_add_1981_27 (.A0(n13550), .B0(n28568), .C0(n2897[31]), 
          .D0(n2831_adj_857), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n30771), .S0(n2996[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_27.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_27.INIT1 = 16'h0000;
    defparam div_9_add_1981_27.INJECT1_0 = "NO";
    defparam div_9_add_1981_27.INJECT1_1 = "NO";
    CCU2C div_13_add_1579_17 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[27]), 
          .D0(n2241), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[28]), 
          .D1(n2240), .CIN(n30936), .COUT(n30937), .S0(n2402[27]), .S1(n2402[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1579_17.INJECT1_0 = "NO";
    defparam div_13_add_1579_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_71 (.A(n2344), .B(n2342), .C(n2341), .D(n2336), 
         .Z(n35620)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_71.init = 16'hfffe;
    LUT4 rem_10_i1857_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[23]), 
         .D(n2740), .Z(n2839)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1857_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_72 (.A(n2348), .B(n28315), .C(n2347), .D(n2349), 
         .Z(n28442)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_72.init = 16'h8000;
    LUT4 i23443_2_lut_3_lut (.A(n69_adj_12), .B(n3), .C(n27382), .Z(duty0_14__N_426[5])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23443_2_lut_3_lut.init = 16'he0e0;
    CCU2C div_9_add_1378_3 (.A0(n13613), .B0(n28526), .C0(n2006_adj_2170[16]), 
          .D0(n335), .A1(n13613), .B1(n28526), .C1(n2006_adj_2170[17]), 
          .D1(n1954_adj_863), .CIN(n30654), .COUT(n30655), .S0(n2105[16]), 
          .S1(n2105[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1378_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1378_3.INJECT1_0 = "NO";
    defparam div_9_add_1378_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1579_15 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[25]), 
          .D0(n2243), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[26]), 
          .D1(n2242), .CIN(n30935), .COUT(n30936), .S0(n2402[25]), .S1(n2402[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1579_15.INJECT1_0 = "NO";
    defparam div_13_add_1579_15.INJECT1_1 = "NO";
    LUT4 i24362_4_lut (.A(n2351), .B(n2350), .C(n28058), .D(n2352), 
         .Z(n28315)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24362_4_lut.init = 16'heccc;
    LUT4 i24108_3_lut (.A(n339), .B(n2353), .C(n2354), .Z(n28058)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24108_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_73 (.A(n36338), .B(n1943_adj_777), .C(n1940_adj_758), 
         .D(n1942_adj_779), .Z(n13613)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_73.init = 16'hfffe;
    LUT4 i1_4_lut_adj_74 (.A(n1944_adj_785), .B(n1941_adj_756), .C(n1945_adj_783), 
         .D(n1946_adj_802), .Z(n36338)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_74.init = 16'hfffe;
    LUT4 i1_4_lut_adj_75 (.A(n1947_adj_800), .B(n28249), .C(n1948_adj_829), 
         .D(n1949_adj_827), .Z(n28526)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_75.init = 16'h8000;
    CCU2C add_26228_13 (.A0(n108), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n105), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30520), 
          .COUT(n30521), .S0(n38[11]), .S1(n38[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_13.INIT0 = 16'h5550;
    defparam add_26228_13.INIT1 = 16'h5550;
    defparam add_26228_13.INJECT1_0 = "NO";
    defparam add_26228_13.INJECT1_1 = "NO";
    LUT4 i24296_4_lut (.A(n1951_adj_833), .B(n1950_adj_835), .C(n27990), 
         .D(n1952_adj_840), .Z(n28249)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24296_4_lut.init = 16'heccc;
    CCU2C div_9_add_1981_25 (.A0(n13550), .B0(n28568), .C0(n2897[29]), 
          .D0(n38230), .A1(n13550), .B1(n28568), .C1(n2897[30]), .D1(n2832), 
          .CIN(n30770), .COUT(n30771), .S0(n2996[29]), .S1(n2996[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_25.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_25.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_25.INJECT1_0 = "NO";
    defparam div_9_add_1981_25.INJECT1_1 = "NO";
    LUT4 i24040_3_lut (.A(n335), .B(n1953_adj_838), .C(n1954_adj_863), 
         .Z(n27990)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24040_3_lut.init = 16'hecec;
    LUT4 i23489_2_lut_rep_328 (.A(n72_adj_13), .B(n3), .Z(n38333)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23489_2_lut_rep_328.init = 16'heeee;
    LUT4 rem_10_i1853_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[27]), 
         .D(n38244), .Z(n2835)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1853_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23444_2_lut_3_lut (.A(n72_adj_13), .B(n3), .C(n27382), .Z(duty0_14__N_426[4])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23444_2_lut_3_lut.init = 16'he0e0;
    CCU2C div_13_add_1579_13 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[23]), 
          .D0(n2245), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[24]), 
          .D1(n2244), .CIN(n30934), .COUT(n30935), .S0(n2402[23]), .S1(n2402[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1579_13.INJECT1_0 = "NO";
    defparam div_13_add_1579_13.INJECT1_1 = "NO";
    CCU2C div_9_add_1378_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n45), .D1(n35[15]), 
          .COUT(n30654), .S1(n2105[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1378_1.INIT0 = 16'h0000;
    defparam div_9_add_1378_1.INIT1 = 16'habef;
    defparam div_9_add_1378_1.INJECT1_0 = "NO";
    defparam div_9_add_1378_1.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_51_i27_2_lut (.A(pwm_cnt[13]), .B(duty3[13]), .Z(n36927)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i27_2_lut.init = 16'h9999;
    CCU2C div_9_add_1311_17 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[31]), 
          .D0(n1841_adj_874), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n30653), .S0(n2006_adj_2170[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1311_17.INIT1 = 16'h0000;
    defparam div_9_add_1311_17.INJECT1_0 = "NO";
    defparam div_9_add_1311_17.INJECT1_1 = "NO";
    LUT4 div_9_i2264_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[18]), 
         .D(n3339_adj_875), .Z(n37)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2264_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1579_11 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[21]), 
          .D0(n2247), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[22]), 
          .D1(n2246), .CIN(n30933), .COUT(n30934), .S0(n2402[21]), .S1(n2402[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1579_11.INJECT1_0 = "NO";
    defparam div_13_add_1579_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1981_23 (.A0(n13550), .B0(n28568), .C0(n2897[27]), 
          .D0(n38231), .A1(n13550), .B1(n28568), .C1(n2897[28]), .D1(n2834_adj_880), 
          .CIN(n30769), .COUT(n30770), .S0(n2996[27]), .S1(n2996[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_23.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_23.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_23.INJECT1_0 = "NO";
    defparam div_9_add_1981_23.INJECT1_1 = "NO";
    CCU2C div_13_add_1579_9 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[19]), 
          .D0(n2249), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[20]), 
          .D1(n2248), .CIN(n30932), .COUT(n30933), .S0(n2402[19]), .S1(n2402[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1579_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1579_9.INJECT1_0 = "NO";
    defparam div_13_add_1579_9.INJECT1_1 = "NO";
    LUT4 rem_10_i1850_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[30]), 
         .D(n2733_adj_884), .Z(n2832_adj_534)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1850_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1981_21 (.A0(n13550), .B0(n28568), .C0(n2897[25]), 
          .D0(n2837_adj_886), .A1(n13550), .B1(n28568), .C1(n2897[26]), 
          .D1(n2836_adj_888), .CIN(n30768), .COUT(n30769), .S0(n2996[25]), 
          .S1(n2996[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_21.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_21.INJECT1_0 = "NO";
    defparam div_9_add_1981_21.INJECT1_1 = "NO";
    LUT4 rem_10_i1860_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[20]), 
         .D(n2743_adj_890), .Z(n2842)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1860_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32202_4_lut (.A(n38374), .B(n36927), .C(n38376), .D(n36891), 
         .Z(n36947)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32202_4_lut.init = 16'hbfbb;
    LUT4 rem_10_i1859_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[21]), 
         .D(n2742_adj_892), .Z(n2841)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1859_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23492_2_lut_rep_329 (.A(n78_adj_14), .B(n3), .Z(n38334)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23492_2_lut_rep_329.init = 16'heeee;
    CCU2C div_9_add_1981_19 (.A0(n13550), .B0(n28568), .C0(n2897[23]), 
          .D0(n2839_adj_665), .A1(n13550), .B1(n28568), .C1(n2897[24]), 
          .D1(n2838), .CIN(n30767), .COUT(n30768), .S0(n2996[23]), .S1(n2996[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_19.INJECT1_0 = "NO";
    defparam div_9_add_1981_19.INJECT1_1 = "NO";
    CCU2C div_13_add_1579_7 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[17]), 
          .D0(n2251), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[18]), 
          .D1(n2250), .CIN(n30931), .COUT(n30932), .S0(n2402[17]), .S1(n2402[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1579_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1579_7.INJECT1_0 = "NO";
    defparam div_13_add_1579_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1981_17 (.A0(n13550), .B0(n28568), .C0(n2897[21]), 
          .D0(n38236), .A1(n13550), .B1(n28568), .C1(n2897[22]), .D1(n2840_adj_899), 
          .CIN(n30766), .COUT(n30767), .S0(n2996[21]), .S1(n2996[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_17.INJECT1_0 = "NO";
    defparam div_9_add_1981_17.INJECT1_1 = "NO";
    CCU2C div_13_add_1579_5 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[15]), 
          .D0(n2253), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[16]), 
          .D1(n2252), .CIN(n30930), .COUT(n30931), .S0(n2402[15]), .S1(n2402[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1579_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1579_5.INJECT1_0 = "NO";
    defparam div_13_add_1579_5.INJECT1_1 = "NO";
    CCU2C div_9_add_1981_15 (.A0(n13550), .B0(n28568), .C0(n2897[19]), 
          .D0(n2843_adj_903), .A1(n13550), .B1(n28568), .C1(n2897[20]), 
          .D1(n2842_adj_764), .CIN(n30765), .COUT(n30766), .S0(n2996[19]), 
          .S1(n2996[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_15.INJECT1_0 = "NO";
    defparam div_9_add_1981_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_1445_15 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[26]), 
          .D0(n2044_adj_905), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[27]), 
          .D1(n38280), .CIN(n30577), .COUT(n30578), .S0(n2204_adj_2172[26]), 
          .S1(n2204_adj_2172[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1445_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1445_15.INJECT1_0 = "NO";
    defparam rem_10_add_1445_15.INJECT1_1 = "NO";
    LUT4 i23451_2_lut_3_lut (.A(n78_adj_14), .B(n3), .C(n27382), .Z(duty0_14__N_426[2])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23451_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_4_lut_adj_76 (.A(n35516), .B(n35514), .C(n2244), .D(n2240), 
         .Z(n13633)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_76.init = 16'hfffe;
    CCU2C add_26228_11 (.A0(n114), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n111), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30519), 
          .COUT(n30520), .S0(n38[9]), .S1(n38[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_11.INIT0 = 16'h5550;
    defparam add_26228_11.INIT1 = 16'h5550;
    defparam add_26228_11.INJECT1_0 = "NO";
    defparam add_26228_11.INJECT1_1 = "NO";
    LUT4 rem_10_i1865_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[15]), 
         .D(n2748_adj_911), .Z(n2847)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1865_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_77 (.A(n2245), .B(n2246), .C(n2239), .D(n2242), 
         .Z(n35516)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_77.init = 16'hfffe;
    LUT4 i1_4_lut_adj_78 (.A(n2243), .B(n2237), .C(n2238), .D(n2241), 
         .Z(n35514)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_78.init = 16'hfffe;
    LUT4 i1_4_lut_adj_79 (.A(n2248), .B(n28317), .C(n2247), .D(n2249), 
         .Z(n28430)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_79.init = 16'h8000;
    CCU2C div_13_add_1579_3 (.A0(n13633), .B0(n28430), .C0(n2303_adj_2171[13]), 
          .D0(n338_adj_913), .A1(n13633), .B1(n28430), .C1(n2303_adj_2171[14]), 
          .D1(n2254), .CIN(n30929), .COUT(n30930), .S0(n2402[13]), .S1(n2402[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1579_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1579_3.INJECT1_0 = "NO";
    defparam div_13_add_1579_3.INJECT1_1 = "NO";
    LUT4 i24364_4_lut (.A(n2251), .B(n2250), .C(n28060), .D(n2252), 
         .Z(n28317)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24364_4_lut.init = 16'heccc;
    LUT4 i23493_2_lut_rep_330 (.A(n81_adj_15), .B(n3), .Z(n38335)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23493_2_lut_rep_330.init = 16'heeee;
    CCU2C div_9_add_1981_13 (.A0(n13550), .B0(n28568), .C0(n2897[17]), 
          .D0(n2845_adj_917), .A1(n13550), .B1(n28568), .C1(n2897[18]), 
          .D1(n2844_adj_919), .CIN(n30764), .COUT(n30765), .S0(n2996[17]), 
          .S1(n2996[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_13.INJECT1_0 = "NO";
    defparam div_9_add_1981_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1579_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n339), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30929), .S1(n2402[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1579_1.INIT0 = 16'h0000;
    defparam div_13_add_1579_1.INIT1 = 16'h555a;
    defparam div_13_add_1579_1.INJECT1_0 = "NO";
    defparam div_13_add_1579_1.INJECT1_1 = "NO";
    LUT4 i24110_3_lut (.A(n338_adj_913), .B(n2253), .C(n2254), .Z(n28060)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24110_3_lut.init = 16'hecec;
    CCU2C add_26228_9 (.A0(n120), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n117), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30518), 
          .COUT(n30519), .S0(n38[7]), .S1(n38[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_9.INIT0 = 16'h5550;
    defparam add_26228_9.INIT1 = 16'h5550;
    defparam add_26228_9.INJECT1_0 = "NO";
    defparam add_26228_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_80 (.A(n2040_adj_844), .B(n35694), .C(n35692), .D(n2045_adj_922), 
         .Z(n13595)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_80.init = 16'hfffe;
    LUT4 i23453_2_lut_3_lut (.A(n81_adj_15), .B(n3), .C(n27382), .Z(duty0_14__N_426[1])) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(54[16] 56[10])
    defparam i23453_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_4_lut_adj_81 (.A(n2041_adj_850), .B(n2044_adj_905), .C(n2046), 
         .D(n2039_adj_845), .Z(n35694)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_81.init = 16'hfffe;
    LUT4 i1_4_lut_adj_82 (.A(n2047_adj_923), .B(n28168), .C(n2048_adj_924), 
         .D(n2049_adj_925), .Z(n28407)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_82.init = 16'h8000;
    LUT4 i24216_4_lut (.A(n2051_adj_926), .B(n2050_adj_927), .C(n27890), 
         .D(n2052_adj_928), .Z(n28168)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24216_4_lut.init = 16'heccc;
    CCU2C div_13_add_1512_19 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[30]), 
          .D0(n2139), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[31]), 
          .D1(n2138), .CIN(n30927), .S0(n2303_adj_2171[30]), .S1(n2303_adj_2171[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1512_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1512_19.INJECT1_0 = "NO";
    defparam div_13_add_1512_19.INJECT1_1 = "NO";
    LUT4 i23941_3_lut (.A(n585), .B(n2053_adj_931), .C(n2054_adj_932), 
         .Z(n27890)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23941_3_lut.init = 16'hecec;
    CCU2C div_9_add_1981_11 (.A0(n13550), .B0(n28568), .C0(n2897[15]), 
          .D0(n2847_adj_934), .A1(n13550), .B1(n28568), .C1(n2897[16]), 
          .D1(n2846_adj_936), .CIN(n30763), .COUT(n30764), .S0(n2996[15]), 
          .S1(n2996[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_11.INJECT1_0 = "NO";
    defparam div_9_add_1981_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_83 (.A(n3132), .B(n3194_adj_2175[27]), .C(n38199), 
         .D(n3240_adj_561), .Z(n35264)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_83.init = 16'hffca;
    LUT4 i1_4_lut_adj_84 (.A(n36208), .B(n36186), .C(n36202), .D(n36196), 
         .Z(n13550)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_84.init = 16'hfffe;
    CCU2C div_9_add_1981_9 (.A0(n13550), .B0(n28568), .C0(n2897[13]), 
          .D0(n2849_adj_939), .A1(n13550), .B1(n28568), .C1(n2897[14]), 
          .D1(n2848), .CIN(n30762), .COUT(n30763), .S0(n2996[13]), .S1(n2996[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1981_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1981_9.INJECT1_0 = "NO";
    defparam div_9_add_1981_9.INJECT1_1 = "NO";
    LUT4 rem_10_i1866_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[14]), 
         .D(n2749_adj_941), .Z(n2848_adj_570)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1866_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1867_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[13]), 
         .D(n2750_adj_943), .Z(n2849)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1867_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1871_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[9]), 
         .D(n2754_adj_945), .Z(n2853)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1871_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_85 (.A(n2840_adj_899), .B(n36204), .C(n36188), .D(n2837_adj_886), 
         .Z(n36208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_85.init = 16'hfffe;
    LUT4 rem_10_i1872_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[8]), 
         .D(n592), .Z(n2854)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1872_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_86 (.A(n2836_adj_888), .B(n2844_adj_919), .C(n2846_adj_936), 
         .D(n2843_adj_903), .Z(n36202)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_86.init = 16'hfffe;
    LUT4 rem_10_i1869_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[11]), 
         .D(n38246), .Z(n2851)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1869_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_87 (.A(n3030), .B(n3095_adj_2176[30]), .C(n38195), 
         .D(n3139_adj_753), .Z(n35342)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_87.init = 16'hffca;
    LUT4 i1_4_lut_adj_88 (.A(n2845_adj_917), .B(n2831_adj_857), .C(n2834_adj_880), 
         .D(n2838), .Z(n36204)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_88.init = 16'hfffe;
    LUT4 i1_4_lut_adj_89 (.A(n2847_adj_934), .B(n28508), .C(n2848), .D(n2849_adj_939), 
         .Z(n28568)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_89.init = 16'h8000;
    LUT4 rem_10_i1868_3_lut_4_lut (.A(n28373), .B(n13626), .C(n2798_adj_2165[12]), 
         .D(n2751_adj_950), .Z(n2850)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1868_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24554_4_lut (.A(n2851_adj_951), .B(n2850_adj_952), .C(n28210), 
         .D(n2852_adj_953), .Z(n28508)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24554_4_lut.init = 16'heccc;
    LUT4 i24258_3_lut (.A(n344), .B(n2853_adj_954), .C(n2854_adj_955), 
         .Z(n28210)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24258_3_lut.init = 16'hecec;
    LUT4 i24602_2_lut_rep_235 (.A(n28554), .B(n13551), .Z(n38240)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24602_2_lut_rep_235.init = 16'heeee;
    LUT4 i1_4_lut_adj_90 (.A(n1841_adj_874), .B(n1844), .C(n1846_adj_956), 
         .D(n1842_adj_957), .Z(n36346)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_90.init = 16'hfffe;
    LUT4 i1_4_lut_adj_91 (.A(n1847_adj_958), .B(n28257), .C(n1848_adj_959), 
         .D(n1849_adj_960), .Z(n28321)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_91.init = 16'h8000;
    LUT4 div_9_i1859_3_lut_rep_231_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[21]), 
         .D(n2742_adj_762), .Z(n38236)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1859_3_lut_rep_231_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1853_3_lut_rep_226_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[27]), 
         .D(n2736_adj_663), .Z(n38231)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1853_3_lut_rep_226_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1311_15 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[29]), 
          .D0(n1843), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[30]), 
          .D1(n1842_adj_957), .CIN(n30652), .COUT(n30653), .S0(n2006_adj_2170[29]), 
          .S1(n2006_adj_2170[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1311_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1311_15.INJECT1_0 = "NO";
    defparam div_9_add_1311_15.INJECT1_1 = "NO";
    LUT4 i24304_4_lut (.A(n1851_adj_963), .B(n1850_adj_964), .C(n28006), 
         .D(n1852), .Z(n28257)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24304_4_lut.init = 16'heccc;
    LUT4 div_9_i1860_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[20]), 
         .D(n2743_adj_966), .Z(n2842_adj_764)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1860_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24056_3_lut (.A(n334), .B(n1853_adj_967), .C(n1854_adj_968), 
         .Z(n28006)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24056_3_lut.init = 16'hecec;
    CCU2C rem_10_add_1445_13 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[24]), 
          .D0(n2046), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[25]), 
          .D1(n2045_adj_922), .CIN(n30576), .COUT(n30577), .S0(n2204_adj_2172[24]), 
          .S1(n2204_adj_2172[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1445_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1445_13.INJECT1_0 = "NO";
    defparam rem_10_add_1445_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1445_11 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[22]), 
          .D0(n2048_adj_924), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[23]), 
          .D1(n2047_adj_923), .CIN(n30575), .COUT(n30576), .S0(n2204_adj_2172[22]), 
          .S1(n2204_adj_2172[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_11.INIT0 = 16'hf1e0;
    defparam rem_10_add_1445_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1445_11.INJECT1_0 = "NO";
    defparam rem_10_add_1445_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1311_13 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[27]), 
          .D0(n1845_adj_974), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[28]), 
          .D1(n1844), .CIN(n30651), .COUT(n30652), .S0(n2006_adj_2170[27]), 
          .S1(n2006_adj_2170[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1311_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1311_13.INJECT1_0 = "NO";
    defparam div_9_add_1311_13.INJECT1_1 = "NO";
    CCU2C add_26228_7 (.A0(n126), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n123), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30517), 
          .COUT(n30518), .S0(n38[5]), .S1(n38[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_7.INIT0 = 16'h5550;
    defparam add_26228_7.INIT1 = 16'h5550;
    defparam add_26228_7.INJECT1_0 = "NO";
    defparam add_26228_7.INJECT1_1 = "NO";
    CCU2C add_26228_5 (.A0(n132), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n129), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30516), 
          .COUT(n30517), .S0(n38[3]), .S1(n38[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_5.INIT0 = 16'h5550;
    defparam add_26228_5.INIT1 = 16'h5550;
    defparam add_26228_5.INJECT1_0 = "NO";
    defparam add_26228_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_92 (.A(n35660), .B(n35658), .C(n2141_adj_983), .D(n2143_adj_984), 
         .Z(n13634)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_92.init = 16'hfffe;
    LUT4 i1_4_lut_adj_93 (.A(n2146_adj_985), .B(n2144_adj_986), .C(n2139), 
         .D(n2138), .Z(n35660)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_93.init = 16'hfffe;
    CCU2C add_26228_3 (.A0(n138), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n135), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30515), 
          .COUT(n30516), .S0(n38[1]), .S1(n38[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_3.INIT0 = 16'h5550;
    defparam add_26228_3.INIT1 = 16'h5550;
    defparam add_26228_3.INJECT1_0 = "NO";
    defparam add_26228_3.INJECT1_1 = "NO";
    LUT4 div_9_i1868_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[12]), 
         .D(n2751_adj_989), .Z(n2850_adj_952)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1868_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_94 (.A(n2142_adj_990), .B(n2145), .C(n2140_adj_991), 
         .Z(n35658)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_3_lut_adj_94.init = 16'hfefe;
    LUT4 i1_4_lut_adj_95 (.A(n2148_adj_992), .B(n28329), .C(n2147_adj_993), 
         .D(n2149_adj_994), .Z(n28412)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_95.init = 16'h8000;
    LUT4 i24376_4_lut (.A(n2151_adj_995), .B(n2150_adj_996), .C(n28070), 
         .D(n2152), .Z(n28329)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24376_4_lut.init = 16'heccc;
    LUT4 div_9_i1852_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[28]), 
         .D(n2735_adj_998), .Z(n2834_adj_880)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1852_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1981_7 (.A0(n13550), .B0(n28568), .C0(n2897[11]), 
          .D0(n2851_adj_951), .A1(n13550), .B1(n28568), .C1(n2897[12]), 
          .D1(n2850_adj_952), .CIN(n30761), .COUT(n30762), .S0(n2996[11]), 
          .S1(n2996[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1981_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1981_7.INJECT1_0 = "NO";
    defparam div_9_add_1981_7.INJECT1_1 = "NO";
    CCU2C add_26228_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n141), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .COUT(n30515));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_26228_1.INIT0 = 16'h0000;
    defparam add_26228_1.INIT1 = 16'haaaf;
    defparam add_26228_1.INJECT1_0 = "NO";
    defparam add_26228_1.INJECT1_1 = "NO";
    LUT4 i24120_3_lut (.A(n337_adj_1001), .B(n2153_adj_1002), .C(n2154_adj_1003), 
         .Z(n28070)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24120_3_lut.init = 16'hecec;
    CCU2C rem_10_add_1445_9 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[20]), 
          .D0(n2050_adj_927), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[21]), 
          .D1(n2049_adj_925), .CIN(n30574), .COUT(n30575), .S0(n2204_adj_2172[20]), 
          .S1(n2204_adj_2172[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1445_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1445_9.INJECT1_0 = "NO";
    defparam rem_10_add_1445_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_17 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[28]), 
          .D0(n2141_adj_983), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[29]), 
          .D1(n2140_adj_991), .CIN(n30926), .COUT(n30927), .S0(n2303_adj_2171[28]), 
          .S1(n2303_adj_2171[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1512_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1512_17.INJECT1_0 = "NO";
    defparam div_13_add_1512_17.INJECT1_1 = "NO";
    CCU2C div_9_add_1311_11 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[25]), 
          .D0(n1847_adj_958), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[26]), 
          .D1(n1846_adj_956), .CIN(n30650), .COUT(n30651), .S0(n2006_adj_2170[25]), 
          .S1(n2006_adj_2170[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1311_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1311_11.INJECT1_0 = "NO";
    defparam div_9_add_1311_11.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_15 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[26]), 
          .D0(n2143_adj_984), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[27]), 
          .D1(n2142_adj_990), .CIN(n30925), .COUT(n30926), .S0(n2303_adj_2171[26]), 
          .S1(n2303_adj_2171[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1512_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1512_15.INJECT1_0 = "NO";
    defparam div_13_add_1512_15.INJECT1_1 = "NO";
    CCU2C div_9_add_1981_5 (.A0(n13550), .B0(n28568), .C0(n2897[9]), .D0(n2853_adj_954), 
          .A1(n13550), .B1(n28568), .C1(n2897[10]), .D1(n2852_adj_953), 
          .CIN(n30760), .COUT(n30761), .S0(n2996[9]), .S1(n2996[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1981_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1981_5.INJECT1_0 = "NO";
    defparam div_9_add_1981_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_96 (.A(n36160), .B(n36178), .C(n36176), .D(n2736_adj_663), 
         .Z(n13551)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_96.init = 16'hfffe;
    CCU2C rem_10_add_1445_7 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[18]), 
          .D0(n2052_adj_928), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[19]), 
          .D1(n2051_adj_926), .CIN(n30573), .COUT(n30574), .S0(n2204_adj_2172[18]), 
          .S1(n2204_adj_2172[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_7.INIT0 = 16'hf1e0;
    defparam rem_10_add_1445_7.INIT1 = 16'h0e1f;
    defparam rem_10_add_1445_7.INJECT1_0 = "NO";
    defparam rem_10_add_1445_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_13 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[24]), 
          .D0(n2145), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[25]), 
          .D1(n2144_adj_986), .CIN(n30924), .COUT(n30925), .S0(n2303_adj_2171[24]), 
          .S1(n2303_adj_2171[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1512_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1512_13.INJECT1_0 = "NO";
    defparam div_13_add_1512_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_97 (.A(n2737_adj_1018), .B(n36174), .C(n36168), 
         .D(n2733_adj_1019), .Z(n36178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_97.init = 16'hfffe;
    CCU2C div_9_add_1981_3 (.A0(n13550), .B0(n28568), .C0(n2897[7]), .D0(n344), 
          .A1(n13550), .B1(n28568), .C1(n2897[8]), .D1(n2854_adj_955), 
          .CIN(n30759), .COUT(n30760), .S0(n2996[7]), .S1(n2996[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1981_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1981_3.INJECT1_0 = "NO";
    defparam div_9_add_1981_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1445_5 (.A0(n13595), .B0(n28407), .C0(n2105_adj_2168[16]), 
          .D0(n2054_adj_932), .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[17]), 
          .D1(n2053_adj_931), .CIN(n30572), .COUT(n30573), .S0(n2204_adj_2172[16]), 
          .S1(n2204_adj_2172[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_5.INIT0 = 16'h0e1f;
    defparam rem_10_add_1445_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1445_5.INJECT1_0 = "NO";
    defparam rem_10_add_1445_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1445_3 (.A0(n12154), .B0(n5), .C0(n48), .D0(n2[14]), 
          .A1(n13595), .B1(n28407), .C1(n2105_adj_2168[15]), .D1(n585), 
          .CIN(n30571), .COUT(n30572), .S0(n2204_adj_2172[14]), .S1(n2204_adj_2172[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_3.INIT0 = 16'h5410;
    defparam rem_10_add_1445_3.INIT1 = 16'hf1e0;
    defparam rem_10_add_1445_3.INJECT1_0 = "NO";
    defparam rem_10_add_1445_3.INJECT1_1 = "NO";
    CCU2C div_9_add_1981_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[6]), .D1(duty0_14__N_426[4]), 
          .COUT(n30759), .S1(n2996[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1981_1.INIT0 = 16'h0000;
    defparam div_9_add_1981_1.INIT1 = 16'h04bf;
    defparam div_9_add_1981_1.INJECT1_0 = "NO";
    defparam div_9_add_1981_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1311_9 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[23]), 
          .D0(n1849_adj_960), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[24]), 
          .D1(n1848_adj_959), .CIN(n30649), .COUT(n30650), .S0(n2006_adj_2170[23]), 
          .S1(n2006_adj_2170[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1311_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1311_9.INJECT1_0 = "NO";
    defparam div_9_add_1311_9.INJECT1_1 = "NO";
    CCU2C div_9_add_1311_7 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[21]), 
          .D0(n1851_adj_963), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[22]), 
          .D1(n1850_adj_964), .CIN(n30648), .COUT(n30649), .S0(n2006_adj_2170[21]), 
          .S1(n2006_adj_2170[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1311_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1311_7.INJECT1_0 = "NO";
    defparam div_9_add_1311_7.INJECT1_1 = "NO";
    LUT4 i24473_2_lut_3_lut_4_lut (.A(n28512), .B(n13602), .C(n33356), 
         .D(n38164), .Z(n60_adj_1030)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam i24473_2_lut_3_lut_4_lut.init = 16'h000e;
    LUT4 div_9_i1861_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[19]), 
         .D(n2744_adj_1032), .Z(n2843_adj_903)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1861_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_98 (.A(n2744_adj_1032), .B(n2742_adj_762), .C(n2745_adj_1033), 
         .D(n2746_adj_1034), .Z(n36176)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_98.init = 16'hfffe;
    LUT4 i1_4_lut_adj_99 (.A(n2743_adj_966), .B(n2735_adj_998), .C(n2739_adj_1035), 
         .D(n2741_adj_1036), .Z(n36174)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_99.init = 16'hfffe;
    LUT4 div_9_i1871_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[9]), 
         .D(n2754_adj_1038), .Z(n2853_adj_954)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1871_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_100 (.A(n2747_adj_1039), .B(n28510), .C(n2748_adj_1040), 
         .D(n2749_adj_1041), .Z(n28554)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_100.init = 16'h8000;
    LUT4 div_9_i1870_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[10]), 
         .D(n2753_adj_1043), .Z(n2852_adj_953)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1870_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1865_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[15]), 
         .D(n2748_adj_1040), .Z(n2847_adj_934)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1865_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_101 (.A(n3031), .B(n3095_adj_2176[29]), .C(n38195), 
         .D(n3143), .Z(n35338)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_101.init = 16'hffca;
    LUT4 i24556_4_lut (.A(n2751_adj_989), .B(n2750_adj_1046), .C(n28214), 
         .D(n2752_adj_1047), .Z(n28510)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24556_4_lut.init = 16'heccc;
    LUT4 i24262_3_lut (.A(n343_adj_677), .B(n2753_adj_1043), .C(n2754_adj_1038), 
         .Z(n28214)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24262_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_102 (.A(n2045_adj_1048), .B(n35716), .C(n35714), 
         .D(n2043_adj_1049), .Z(n13635)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_102.init = 16'hfffe;
    LUT4 div_9_i1851_3_lut_rep_225_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[29]), 
         .D(n2734_adj_650), .Z(n38230)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1851_3_lut_rep_225_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_103 (.A(n2044_adj_1050), .B(n2040_adj_1051), .C(n2046_adj_1052), 
         .D(n2042_adj_1053), .Z(n35716)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_103.init = 16'hfffe;
    LUT4 div_9_i1867_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[13]), 
         .D(n2750_adj_1046), .Z(n2849_adj_939)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1867_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_104 (.A(n3033_adj_1055), .B(n3095_adj_2176[27]), 
         .C(n38195), .D(n3137_adj_674), .Z(n35348)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_104.init = 16'hffca;
    LUT4 div_9_i1862_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[18]), 
         .D(n2745_adj_1033), .Z(n2844_adj_919)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1862_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_105 (.A(n2048_adj_1058), .B(n28337), .C(n2047_adj_1059), 
         .D(n2049_adj_1060), .Z(n28401)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_105.init = 16'h8000;
    LUT4 i24384_4_lut (.A(n2051_adj_1061), .B(n2050_adj_1062), .C(n27972), 
         .D(n2052_adj_1063), .Z(n28337)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24384_4_lut.init = 16'heccc;
    LUT4 i24022_3_lut (.A(n336_adj_1064), .B(n2053_adj_1065), .C(n2054_adj_1066), 
         .Z(n27972)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24022_3_lut.init = 16'hecec;
    LUT4 i26579_4_lut (.A(n38305), .B(n35960), .C(n1709_adj_2160[30]), 
         .D(n1709_adj_2160[28]), .Z(n13653)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i26579_4_lut.init = 16'haaa8;
    LUT4 div_9_i1869_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[11]), 
         .D(n2752_adj_1047), .Z(n2851_adj_951)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1869_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_106 (.A(n1709_adj_2160[29]), .B(n1709_adj_2160[31]), 
         .C(n1709_adj_2160[27]), .Z(n35960)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_3_lut_adj_106.init = 16'hfefe;
    LUT4 div_9_i1872_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[8]), 
         .D(n343_adj_677), .Z(n2854_adj_955)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1872_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_107 (.A(n35834), .B(n1750_adj_1073), .C(n1709_adj_2160[26]), 
         .D(n34329), .Z(n28287)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_107.init = 16'ha080;
    LUT4 i1_4_lut_adj_108 (.A(n35830), .B(n1709_adj_2160[20]), .C(n333), 
         .D(n1754_adj_1076), .Z(n34329)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_108.init = 16'ha888;
    CCU2C div_9_add_1311_5 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[19]), 
          .D0(n1853_adj_967), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[20]), 
          .D1(n1852), .CIN(n30647), .COUT(n30648), .S0(n2006_adj_2170[19]), 
          .S1(n2006_adj_2170[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1311_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1311_5.INJECT1_0 = "NO";
    defparam div_9_add_1311_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(n1709_adj_2160[22]), .B(n1709_adj_2160[21]), .Z(n35830)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 div_9_i1854_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[26]), 
         .D(n2737_adj_1018), .Z(n2836_adj_888)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1854_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_52_i27_2_lut (.A(pwm_cnt[13]), .B(duty2[13]), .Z(n36870)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i27_2_lut.init = 16'h9999;
    LUT4 i24566_2_lut_rep_190 (.A(n28518), .B(n13617), .Z(n38195)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24566_2_lut_rep_190.init = 16'heeee;
    LUT4 div_9_i1857_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[23]), 
         .D(n38245), .Z(n2839_adj_665)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1857_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1914_25 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[30]), 
          .D0(n2733_adj_1019), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[31]), 
          .D1(n38243), .CIN(n30757), .S0(n2897[30]), .S1(n2897[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_25.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_25.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_25.INJECT1_0 = "NO";
    defparam div_9_add_1914_25.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_23 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[28]), 
          .D0(n2735_adj_998), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[29]), 
          .D1(n2734_adj_650), .CIN(n30756), .COUT(n30757), .S0(n2897[28]), 
          .S1(n2897[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_23.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_23.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_23.INJECT1_0 = "NO";
    defparam div_9_add_1914_23.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_21 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[26]), 
          .D0(n2737_adj_1018), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[27]), 
          .D1(n2736_adj_663), .CIN(n30755), .COUT(n30756), .S0(n2897[26]), 
          .S1(n2897[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_21.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_21.INJECT1_0 = "NO";
    defparam div_9_add_1914_21.INJECT1_1 = "NO";
    CCU2C div_9_add_1311_3 (.A0(n38289), .B0(n28321), .C0(n1907_adj_2173[17]), 
          .D0(n334), .A1(n38289), .B1(n28321), .C1(n1907_adj_2173[18]), 
          .D1(n1854_adj_968), .CIN(n30646), .COUT(n30647), .S0(n2006_adj_2170[17]), 
          .S1(n2006_adj_2170[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1311_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1311_3.INJECT1_0 = "NO";
    defparam div_9_add_1311_3.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_19 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[24]), 
          .D0(n2739_adj_1035), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[25]), 
          .D1(n2738_adj_1089), .CIN(n30754), .COUT(n30755), .S0(n2897[24]), 
          .S1(n2897[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_19.INJECT1_0 = "NO";
    defparam div_9_add_1914_19.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_11 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[22]), 
          .D0(n2147_adj_993), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[23]), 
          .D1(n2146_adj_985), .CIN(n30923), .COUT(n30924), .S0(n2303_adj_2171[22]), 
          .S1(n2303_adj_2171[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1512_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1512_11.INJECT1_0 = "NO";
    defparam div_13_add_1512_11.INJECT1_1 = "NO";
    LUT4 n3397_bdd_4_lut_32259 (.A(n3392_adj_2177[27]), .B(n3392_adj_2177[19]), 
         .C(n3392_adj_2177[29]), .D(n3392_adj_2177[20]), .Z(n37486)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3397_bdd_4_lut_32259.init = 16'hfffe;
    LUT4 div_9_i1863_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[17]), 
         .D(n2746_adj_1034), .Z(n2845_adj_917)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1863_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2054_3_lut_rep_189_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[27]), 
         .D(n3033_adj_1055), .Z(n38194)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2054_3_lut_rep_189_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1864_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[16]), 
         .D(n2747_adj_1039), .Z(n2846_adj_936)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1864_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2052_3_lut_rep_188_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[29]), 
         .D(n3031), .Z(n38193)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2052_3_lut_rep_188_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1849_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[31]), 
         .D(n38243), .Z(n2831_adj_857)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1849_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2411_3_lut_4_lut (.A(n28554), .B(n13551), .C(n38307), 
         .D(n4540[7]), .Z(n89[7])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_9_i2411_3_lut_4_lut.init = 16'hfe0e;
    LUT4 div_9_i1858_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[22]), 
         .D(n2741_adj_1036), .Z(n2840_adj_899)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1858_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32204_4_lut (.A(n38370), .B(n36870), .C(n38372), .D(n36834), 
         .Z(n36943)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32204_4_lut.init = 16'hbfbb;
    LUT4 div_9_i1855_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[25]), 
         .D(n2738_adj_1089), .Z(n2837_adj_886)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1855_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1512_9 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[20]), 
          .D0(n2149_adj_994), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[21]), 
          .D1(n2148_adj_992), .CIN(n30922), .COUT(n30923), .S0(n2303_adj_2171[20]), 
          .S1(n2303_adj_2171[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1512_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1512_9.INJECT1_0 = "NO";
    defparam div_13_add_1512_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_7 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[18]), 
          .D0(n2151_adj_995), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[19]), 
          .D1(n2150_adj_996), .CIN(n30921), .COUT(n30922), .S0(n2303_adj_2171[18]), 
          .S1(n2303_adj_2171[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1512_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1512_7.INJECT1_0 = "NO";
    defparam div_13_add_1512_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_5 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[16]), 
          .D0(n2153_adj_1002), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[17]), 
          .D1(n2152), .CIN(n30920), .COUT(n30921), .S0(n2303_adj_2171[16]), 
          .S1(n2303_adj_2171[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1512_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1512_5.INJECT1_0 = "NO";
    defparam div_13_add_1512_5.INJECT1_1 = "NO";
    CCU2C div_13_add_1512_3 (.A0(n13634), .B0(n28412), .C0(n2204_adj_2174[14]), 
          .D0(n337_adj_1001), .A1(n13634), .B1(n28412), .C1(n2204_adj_2174[15]), 
          .D1(n2154_adj_1003), .CIN(n30919), .COUT(n30920), .S0(n2303_adj_2171[14]), 
          .S1(n2303_adj_2171[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1512_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1512_3.INJECT1_0 = "NO";
    defparam div_13_add_1512_3.INJECT1_1 = "NO";
    LUT4 div_9_i1850_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[30]), 
         .D(n2733_adj_1019), .Z(n2832)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1850_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1512_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n338_adj_913), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30919), .S1(n2303_adj_2171[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1512_1.INIT0 = 16'h0000;
    defparam div_13_add_1512_1.INIT1 = 16'h555a;
    defparam div_13_add_1512_1.INJECT1_0 = "NO";
    defparam div_13_add_1512_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1445_19 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[31]), 
          .D0(n38273), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30918), .S0(n2204_adj_2174[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1445_19.INIT1 = 16'h0000;
    defparam div_13_add_1445_19.INJECT1_0 = "NO";
    defparam div_13_add_1445_19.INJECT1_1 = "NO";
    CCU2C div_13_add_1445_17 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[29]), 
          .D0(n2041_adj_1109), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[30]), 
          .D1(n2040_adj_1051), .CIN(n30917), .COUT(n30918), .S0(n2204_adj_2174[29]), 
          .S1(n2204_adj_2174[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1445_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1445_17.INJECT1_0 = "NO";
    defparam div_13_add_1445_17.INJECT1_1 = "NO";
    CCU2C div_9_add_1311_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n42), .D1(n35[16]), 
          .COUT(n30646), .S1(n2006_adj_2170[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1311_1.INIT0 = 16'h0000;
    defparam div_9_add_1311_1.INIT1 = 16'habef;
    defparam div_9_add_1311_1.INJECT1_0 = "NO";
    defparam div_9_add_1311_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_17 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[22]), 
          .D0(n2741_adj_1036), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[23]), 
          .D1(n38245), .CIN(n30753), .COUT(n30754), .S0(n2897[22]), 
          .S1(n2897[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_17.INJECT1_0 = "NO";
    defparam div_9_add_1914_17.INJECT1_1 = "NO";
    LUT4 div_9_i2272_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[10]), 
         .D(n3347_adj_1112), .Z(n21_adj_1113)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2272_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2266_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[16]), 
         .D(n3341_adj_1114), .Z(n33)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2266_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2061_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[20]), 
         .D(n3040_adj_1116), .Z(n3139_adj_753)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2061_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1445_15 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[27]), 
          .D0(n2043_adj_1049), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[28]), 
          .D1(n2042_adj_1053), .CIN(n30916), .COUT(n30917), .S0(n2204_adj_2174[27]), 
          .S1(n2204_adj_2174[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1445_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1445_15.INJECT1_0 = "NO";
    defparam div_13_add_1445_15.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_109 (.A(n35706), .B(n1945_adj_1119), .C(n1940_adj_1120), 
         .D(n1942_adj_1121), .Z(n13636)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_109.init = 16'hfffe;
    LUT4 div_9_i1866_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[14]), 
         .D(n2749_adj_1041), .Z(n2848)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1866_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1856_3_lut_4_lut (.A(n28554), .B(n13551), .C(n2798_adj_2166[24]), 
         .D(n2739_adj_1035), .Z(n2838)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1856_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1445_13 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[25]), 
          .D0(n2045_adj_1048), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[26]), 
          .D1(n2044_adj_1050), .CIN(n30915), .COUT(n30916), .S0(n2204_adj_2174[25]), 
          .S1(n2204_adj_2174[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1445_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1445_13.INJECT1_0 = "NO";
    defparam div_13_add_1445_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_110 (.A(n1944_adj_1125), .B(n1941_adj_1126), .C(n1943_adj_1127), 
         .D(n1946_adj_1128), .Z(n35706)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_110.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_111 (.A(n2534), .B(n2600[31]), .C(n38249), 
         .D(n2634), .Z(n35074)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_111.init = 16'hffca;
    FD1S3IX pwm_cnt_1138__i14 (.D(n50[14]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i14.GSR = "ENABLED";
    CCU2C div_13_add_1445_11 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[23]), 
          .D0(n2047_adj_1059), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[24]), 
          .D1(n2046_adj_1052), .CIN(n30914), .COUT(n30915), .S0(n2204_adj_2174[23]), 
          .S1(n2204_adj_2174[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1445_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1445_11.INJECT1_0 = "NO";
    defparam div_13_add_1445_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_112 (.A(n1948_adj_1132), .B(n28343), .C(n1947_adj_1133), 
         .D(n1949_adj_1134), .Z(n28389)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_112.init = 16'h8000;
    CCU2C div_9_add_1244_15 (.A0(n13653), .B0(n28287), .C0(n1808_adj_2179[30]), 
          .D0(n1743), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[31]), 
          .D1(n1742), .CIN(n30644), .S0(n1907_adj_2173[30]), .S1(n1907_adj_2173[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1244_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1244_15.INJECT1_0 = "NO";
    defparam div_9_add_1244_15.INJECT1_1 = "NO";
    CCU2C div_9_add_1244_13 (.A0(n13653), .B0(n28287), .C0(n1808_adj_2179[28]), 
          .D0(n1745), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[29]), 
          .D1(n1744_adj_520), .CIN(n30643), .COUT(n30644), .S0(n1907_adj_2173[28]), 
          .S1(n1907_adj_2173[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1244_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1244_13.INJECT1_0 = "NO";
    defparam div_9_add_1244_13.INJECT1_1 = "NO";
    LUT4 div_13_i2076_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[5]), 
         .D(n346_adj_1140), .Z(n3154_adj_656)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2076_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1914_15 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[20]), 
          .D0(n2743_adj_966), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[21]), 
          .D1(n2742_adj_762), .CIN(n30752), .COUT(n30753), .S0(n2897[20]), 
          .S1(n2897[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_15.INJECT1_0 = "NO";
    defparam div_9_add_1914_15.INJECT1_1 = "NO";
    CCU2C div_13_add_1445_9 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[21]), 
          .D0(n2049_adj_1060), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[22]), 
          .D1(n2048_adj_1058), .CIN(n30913), .COUT(n30914), .S0(n2204_adj_2174[21]), 
          .S1(n2204_adj_2174[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1445_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1445_9.INJECT1_0 = "NO";
    defparam div_13_add_1445_9.INJECT1_1 = "NO";
    LUT4 i24390_4_lut (.A(n1951_adj_1143), .B(n1950_adj_1144), .C(n28080), 
         .D(n1952_adj_1145), .Z(n28343)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24390_4_lut.init = 16'heccc;
    LUT4 i1_2_lut_4_lut_adj_113 (.A(n2635_adj_1146), .B(n2699_adj_2180[29]), 
         .C(n38248), .D(n2739_adj_816), .Z(n35410)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_113.init = 16'hffca;
    CCU2C div_13_add_1445_7 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[19]), 
          .D0(n2051_adj_1061), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[20]), 
          .D1(n2050_adj_1062), .CIN(n30912), .COUT(n30913), .S0(n2204_adj_2174[19]), 
          .S1(n2204_adj_2174[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1445_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1445_7.INJECT1_0 = "NO";
    defparam div_13_add_1445_7.INJECT1_1 = "NO";
    LUT4 i24129_3_lut (.A(n335_adj_1150), .B(n1953_adj_1151), .C(n1954_adj_1152), 
         .Z(n28080)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24129_3_lut.init = 16'hecec;
    LUT4 i1_3_lut_adj_114 (.A(n27382), .B(n3), .C(n42), .Z(duty0_14__N_426[14])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_114.init = 16'h2020;
    CCU2C div_9_add_1914_13 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[18]), 
          .D0(n2745_adj_1033), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[19]), 
          .D1(n2744_adj_1032), .CIN(n30751), .COUT(n30752), .S0(n2897[18]), 
          .S1(n2897[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_13.INJECT1_0 = "NO";
    defparam div_9_add_1914_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_115 (.A(n36232), .B(n36226), .C(n2635_adj_1153), 
         .D(n2636_adj_1154), .Z(n13552)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_115.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_116 (.A(n2633), .B(n2699_adj_2181[31]), .C(n38247), 
         .D(n2738_adj_1089), .Z(n36160)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_116.init = 16'hffca;
    LUT4 i1_4_lut_adj_117 (.A(n2641_adj_1156), .B(n36228), .C(n36220), 
         .D(n2646_adj_1157), .Z(n36232)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_117.init = 16'hfffe;
    CCU2C div_13_add_1445_5 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[17]), 
          .D0(n2053_adj_1065), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[18]), 
          .D1(n2052_adj_1063), .CIN(n30911), .COUT(n30912), .S0(n2204_adj_2174[17]), 
          .S1(n2204_adj_2174[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1445_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1445_5.INJECT1_0 = "NO";
    defparam div_13_add_1445_5.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_11 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[16]), 
          .D0(n2747_adj_1039), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[17]), 
          .D1(n2746_adj_1034), .CIN(n30750), .COUT(n30751), .S0(n2897[16]), 
          .S1(n2897[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_11.INJECT1_0 = "NO";
    defparam div_9_add_1914_11.INJECT1_1 = "NO";
    CCU2C div_13_add_1445_3 (.A0(n13635), .B0(n28401), .C0(n2105_adj_2178[15]), 
          .D0(n336_adj_1064), .A1(n13635), .B1(n28401), .C1(n2105_adj_2178[16]), 
          .D1(n2054_adj_1066), .CIN(n30910), .COUT(n30911), .S0(n2204_adj_2174[15]), 
          .S1(n2204_adj_2174[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1445_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1445_3.INJECT1_0 = "NO";
    defparam div_13_add_1445_3.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_9 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[14]), 
          .D0(n2749_adj_1041), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[15]), 
          .D1(n2748_adj_1040), .CIN(n30749), .COUT(n30750), .S0(n2897[14]), 
          .S1(n2897[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1914_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1914_9.INJECT1_0 = "NO";
    defparam div_9_add_1914_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_118 (.A(n2640_adj_1162), .B(n2634_adj_1163), .C(n2639_adj_1164), 
         .D(n2638_adj_1165), .Z(n36226)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_118.init = 16'hfffe;
    CCU2C div_9_add_1914_7 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[12]), 
          .D0(n2751_adj_989), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[13]), 
          .D1(n2750_adj_1046), .CIN(n30748), .COUT(n30749), .S0(n2897[12]), 
          .S1(n2897[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1914_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1914_7.INJECT1_0 = "NO";
    defparam div_9_add_1914_7.INJECT1_1 = "NO";
    CCU2C rem_10_add_1445_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n51), .D1(n2[13]), 
          .COUT(n30571));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1445_1.INIT0 = 16'h000F;
    defparam rem_10_add_1445_1.INIT1 = 16'habef;
    defparam rem_10_add_1445_1.INJECT1_0 = "NO";
    defparam rem_10_add_1445_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_119 (.A(n2633), .B(n2637_adj_1166), .C(n2643_adj_1167), 
         .D(n2644_adj_1168), .Z(n36228)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_119.init = 16'hfffe;
    LUT4 i1_4_lut_adj_120 (.A(n2647_adj_1169), .B(n28514), .C(n2648_adj_1170), 
         .D(n2649_adj_1171), .Z(n28544)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_120.init = 16'h8000;
    LUT4 i24560_4_lut (.A(n2651_adj_1172), .B(n2650_adj_1173), .C(n28218), 
         .D(n2652_adj_1174), .Z(n28514)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24560_4_lut.init = 16'heccc;
    LUT4 div_13_i2057_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[24]), 
         .D(n3036_adj_1176), .Z(n3135_adj_687)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2057_3_lut_4_lut.init = 16'hf1e0;
    PFUMX pwm_cnt_14__I_0_52_i28 (.BLUT(n12_adj_1177), .ALUT(n26_adj_1178), 
          .C0(n36943), .Z(n28_adj_1179)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    CCU2C div_13_add_1445_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n337_adj_1001), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30910), .S1(n2204_adj_2174[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1445_1.INIT0 = 16'h0000;
    defparam div_13_add_1445_1.INIT1 = 16'h555a;
    defparam div_13_add_1445_1.INJECT1_0 = "NO";
    defparam div_13_add_1445_1.INJECT1_1 = "NO";
    LUT4 div_13_i2071_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[10]), 
         .D(n3050_adj_1181), .Z(n3149_adj_694)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2071_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2074_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[7]), 
         .D(n3053_adj_1183), .Z(n3152_adj_671)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2074_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24266_3_lut (.A(n342_adj_1184), .B(n2653_adj_1185), .C(n2654_adj_1186), 
         .Z(n28218)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24266_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_121 (.A(n1841_adj_1187), .B(n1844_adj_1188), .C(n1843_adj_1189), 
         .D(n1842_adj_1190), .Z(n35726)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_121.init = 16'hfffe;
    LUT4 i1_4_lut_adj_122 (.A(n1848_adj_1191), .B(n28351), .C(n1847_adj_1192), 
         .D(n1849_adj_1193), .Z(n28377)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_122.init = 16'h8000;
    LUT4 div_13_i2051_3_lut_rep_187_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[30]), 
         .D(n3030), .Z(n38192)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2051_3_lut_rep_187_4_lut.init = 16'hf1e0;
    LUT4 i24398_4_lut (.A(n1851_adj_1194), .B(n1850_adj_1195), .C(n28086), 
         .D(n1852_adj_1196), .Z(n28351)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24398_4_lut.init = 16'heccc;
    CCU2C div_13_add_1378_17 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[30]), 
          .D0(n1941_adj_1126), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[31]), 
          .D1(n1940_adj_1120), .CIN(n30908), .S0(n2105_adj_2178[30]), 
          .S1(n2105_adj_2178[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1378_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1378_17.INJECT1_0 = "NO";
    defparam div_13_add_1378_17.INJECT1_1 = "NO";
    LUT4 i24135_3_lut (.A(n334_adj_1199), .B(n1853_adj_1200), .C(n1854_adj_1201), 
         .Z(n28086)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24135_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_4_lut_adj_123 (.A(n2637_adj_1202), .B(n2699_adj_2180[27]), 
         .C(n38248), .D(n2744_adj_822), .Z(n35402)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_123.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_124 (.A(n2641_adj_1156), .B(n2699_adj_2181[23]), 
         .C(n38247), .D(n2734_adj_650), .Z(n36168)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_124.init = 16'hffca;
    LUT4 pwm_cnt_14__I_0_53_i27_2_lut (.A(pwm_cnt[13]), .B(duty1[13]), .Z(n36813)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i27_2_lut.init = 16'h9999;
    CCU2C div_9_add_1244_11 (.A0(n13653), .B0(n28287), .C0(n1808_adj_2179[26]), 
          .D0(n1747_adj_1206), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[27]), 
          .D1(n1746_adj_1208), .CIN(n30642), .COUT(n30643), .S0(n1907_adj_2173[26]), 
          .S1(n1907_adj_2173[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1244_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1244_11.INJECT1_0 = "NO";
    defparam div_9_add_1244_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_5 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[10]), 
          .D0(n2753_adj_1043), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[11]), 
          .D1(n2752_adj_1047), .CIN(n30747), .COUT(n30748), .S0(n2897[10]), 
          .S1(n2897[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1914_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1914_5.INJECT1_0 = "NO";
    defparam div_9_add_1914_5.INJECT1_1 = "NO";
    LUT4 n3410_bdd_4_lut (.A(n3343_adj_1209), .B(n3341_adj_604), .C(n3347_adj_1210), 
         .D(n3339_adj_565), .Z(n37505)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3410_bdd_4_lut.init = 16'hfffe;
    CCU2C div_9_add_1914_3 (.A0(n13551), .B0(n28554), .C0(n2798_adj_2166[8]), 
          .D0(n343_adj_677), .A1(n13551), .B1(n28554), .C1(n2798_adj_2166[9]), 
          .D1(n2754_adj_1038), .CIN(n30746), .COUT(n30747), .S0(n2897[8]), 
          .S1(n2897[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1914_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1914_3.INJECT1_0 = "NO";
    defparam div_9_add_1914_3.INJECT1_1 = "NO";
    CCU2C div_9_add_1244_9 (.A0(n13653), .B0(n28287), .C0(n1808_adj_2179[24]), 
          .D0(n1749_adj_1212), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[25]), 
          .D1(n38297), .CIN(n30641), .COUT(n30642), .S0(n1907_adj_2173[24]), 
          .S1(n1907_adj_2173[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1244_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1244_9.INJECT1_0 = "NO";
    defparam div_9_add_1244_9.INJECT1_1 = "NO";
    CCU2C div_9_add_1914_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[7]), .D1(duty0_14__N_426[5]), 
          .COUT(n30746), .S1(n2897[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1914_1.INIT0 = 16'h0000;
    defparam div_9_add_1914_1.INIT1 = 16'h04bf;
    defparam div_9_add_1914_1.INJECT1_0 = "NO";
    defparam div_9_add_1914_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_125 (.A(n2653_adj_1214), .B(n2699_adj_2180[11]), 
         .C(n38248), .D(n2751_adj_950), .Z(n34654)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_125.init = 16'hca00;
    LUT4 i24594_2_lut_rep_242 (.A(n28544), .B(n13552), .Z(n38247)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24594_2_lut_rep_242.init = 16'heeee;
    LUT4 div_13_i2066_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[15]), 
         .D(n3045_adj_1217), .Z(n3144_adj_691)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2066_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1378_15 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[28]), 
          .D0(n1943_adj_1127), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[29]), 
          .D1(n1942_adj_1121), .CIN(n30907), .COUT(n30908), .S0(n2105_adj_2178[28]), 
          .S1(n2105_adj_2178[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1378_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1378_15.INJECT1_0 = "NO";
    defparam div_13_add_1378_15.INJECT1_1 = "NO";
    CCU2C div_13_add_1378_13 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[26]), 
          .D0(n1945_adj_1119), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[27]), 
          .D1(n1944_adj_1125), .CIN(n30906), .COUT(n30907), .S0(n2105_adj_2178[26]), 
          .S1(n2105_adj_2178[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1378_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1378_13.INJECT1_0 = "NO";
    defparam div_13_add_1378_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1378_11 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[24]), 
          .D0(n1947_adj_1133), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[25]), 
          .D1(n1946_adj_1128), .CIN(n30905), .COUT(n30906), .S0(n2105_adj_2178[24]), 
          .S1(n2105_adj_2178[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1378_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1378_11.INJECT1_0 = "NO";
    defparam div_13_add_1378_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1847_25 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[31]), 
          .D0(n2633), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30745), .S0(n2798_adj_2166[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_25.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_25.INIT1 = 16'h0000;
    defparam div_9_add_1847_25.INJECT1_0 = "NO";
    defparam div_9_add_1847_25.INJECT1_1 = "NO";
    CCU2C div_9_add_1847_23 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[29]), 
          .D0(n2635_adj_1153), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[30]), 
          .D1(n2634_adj_1163), .CIN(n30744), .COUT(n30745), .S0(n2798_adj_2166[29]), 
          .S1(n2798_adj_2166[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_23.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_23.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_23.INJECT1_0 = "NO";
    defparam div_9_add_1847_23.INJECT1_1 = "NO";
    LUT4 div_9_i1790_3_lut_rep_240_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[23]), 
         .D(n2641_adj_1156), .Z(n38245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1790_3_lut_rep_240_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2059_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[22]), 
         .D(n3038_adj_1227), .Z(n3137_adj_674)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2059_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32206_4_lut (.A(n38366), .B(n36813), .C(n38368), .D(n36777), 
         .Z(n36939)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i32206_4_lut.init = 16'hbfbb;
    CCU2C div_9_add_1244_7 (.A0(n13653), .B0(n28287), .C0(n1808_adj_2179[22]), 
          .D0(n1751_adj_1229), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[23]), 
          .D1(n1750_adj_1073), .CIN(n30640), .COUT(n30641), .S0(n1907_adj_2173[22]), 
          .S1(n1907_adj_2173[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1244_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1244_7.INJECT1_0 = "NO";
    defparam div_9_add_1244_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1378_9 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[22]), 
          .D0(n1949_adj_1134), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[23]), 
          .D1(n1948_adj_1132), .CIN(n30904), .COUT(n30905), .S0(n2105_adj_2178[22]), 
          .S1(n2105_adj_2178[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1378_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1378_9.INJECT1_0 = "NO";
    defparam div_13_add_1378_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_126 (.A(n36308), .B(n36302), .C(n2545_adj_1233), 
         .D(n2546_adj_1234), .Z(n13553)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_126.init = 16'hfffe;
    LUT4 i1_4_lut_adj_127 (.A(n2539_adj_1235), .B(n36304), .C(n2537_adj_1236), 
         .D(n2536_adj_1237), .Z(n36308)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_127.init = 16'hfffe;
    LUT4 i8143_2_lut (.A(n3), .B(n27382), .Z(n12154)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i8143_2_lut.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_128 (.A(n2540_adj_1238), .B(n2544_adj_1239), .C(n2541_adj_1240), 
         .D(n2542_adj_1241), .Z(n36302)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_128.init = 16'hfffe;
    CCU2C div_13_add_1378_7 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[20]), 
          .D0(n1951_adj_1143), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[21]), 
          .D1(n1950_adj_1144), .CIN(n30903), .COUT(n30904), .S0(n2105_adj_2178[20]), 
          .S1(n2105_adj_2178[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1378_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1378_7.INJECT1_0 = "NO";
    defparam div_13_add_1378_7.INJECT1_1 = "NO";
    LUT4 div_9_i1800_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[13]), 
         .D(n2651_adj_1172), .Z(n2750_adj_1046)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1800_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_129 (.A(n2538_adj_1245), .B(n2535_adj_1246), .C(n2543_adj_1247), 
         .D(n2534_adj_1248), .Z(n36304)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_129.init = 16'hfffe;
    LUT4 i1_4_lut_adj_130 (.A(n2547_adj_1249), .B(n28226), .C(n2548_adj_1250), 
         .D(n2549_adj_1251), .Z(n28331)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_130.init = 16'h8000;
    CCU2C div_9_add_1847_21 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[27]), 
          .D0(n2637_adj_1166), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[28]), 
          .D1(n2636_adj_1154), .CIN(n30743), .COUT(n30744), .S0(n2798_adj_2166[27]), 
          .S1(n2798_adj_2166[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_21.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_21.INJECT1_0 = "NO";
    defparam div_9_add_1847_21.INJECT1_1 = "NO";
    CCU2C div_13_add_1378_5 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[18]), 
          .D0(n1953_adj_1151), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[19]), 
          .D1(n1952_adj_1145), .CIN(n30902), .COUT(n30903), .S0(n2105_adj_2178[18]), 
          .S1(n2105_adj_2178[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1378_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1378_5.INJECT1_0 = "NO";
    defparam div_13_add_1378_5.INJECT1_1 = "NO";
    LUT4 div_9_i1801_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[12]), 
         .D(n2652_adj_1174), .Z(n2751_adj_989)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1801_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1847_19 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[25]), 
          .D0(n2639_adj_1164), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[26]), 
          .D1(n2638_adj_1165), .CIN(n30742), .COUT(n30743), .S0(n2798_adj_2166[25]), 
          .S1(n2798_adj_2166[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_19.INJECT1_0 = "NO";
    defparam div_9_add_1847_19.INJECT1_1 = "NO";
    LUT4 i24274_4_lut (.A(n2551_adj_1259), .B(n2550_adj_1260), .C(n27956), 
         .D(n2552_adj_1261), .Z(n28226)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24274_4_lut.init = 16'heccc;
    CCU2C div_13_add_1378_3 (.A0(n13636), .B0(n28389), .C0(n2006_adj_2182[16]), 
          .D0(n335_adj_1150), .A1(n13636), .B1(n28389), .C1(n2006_adj_2182[17]), 
          .D1(n1954_adj_1152), .CIN(n30901), .COUT(n30902), .S0(n2105_adj_2178[16]), 
          .S1(n2105_adj_2178[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1378_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1378_3.INJECT1_0 = "NO";
    defparam div_13_add_1378_3.INJECT1_1 = "NO";
    LUT4 div_13_i2075_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[6]), 
         .D(n3054_adj_1265), .Z(n3153_adj_717)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2075_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1847_17 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[23]), 
          .D0(n2641_adj_1156), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[24]), 
          .D1(n2640_adj_1162), .CIN(n30741), .COUT(n30742), .S0(n2798_adj_2166[23]), 
          .S1(n2798_adj_2166[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_17.INJECT1_0 = "NO";
    defparam div_9_add_1847_17.INJECT1_1 = "NO";
    CCU2C div_13_add_1378_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n336_adj_1064), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30901), .S1(n2105_adj_2178[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1378_1.INIT0 = 16'h0000;
    defparam div_13_add_1378_1.INIT1 = 16'h555a;
    defparam div_13_add_1378_1.INJECT1_0 = "NO";
    defparam div_13_add_1378_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1244_5 (.A0(n13653), .B0(n28287), .C0(n1808_adj_2179[20]), 
          .D0(n1753_adj_1268), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[21]), 
          .D1(n1752_adj_1270), .CIN(n30639), .COUT(n30640), .S0(n1907_adj_2173[20]), 
          .S1(n1907_adj_2173[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1244_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1244_5.INJECT1_0 = "NO";
    defparam div_9_add_1244_5.INJECT1_1 = "NO";
    CCU2C div_13_add_1311_17 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[31]), 
          .D0(n1841_adj_1187), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n30900), .S0(n2006_adj_2182[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1311_17.INIT1 = 16'h0000;
    defparam div_13_add_1311_17.INJECT1_0 = "NO";
    defparam div_13_add_1311_17.INJECT1_1 = "NO";
    LUT4 div_9_i1787_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[26]), 
         .D(n2638_adj_1165), .Z(n2737_adj_1018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1787_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10827_3_lut_4_lut (.A(n28512), .B(n13602), .C(n38307), .D(n4540[1]), 
         .Z(n1)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i10827_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i24006_3_lut (.A(n341), .B(n2553_adj_1272), .C(n2554_adj_1273), 
         .Z(n27956)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24006_3_lut.init = 16'hecec;
    LUT4 div_9_i1802_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[11]), 
         .D(n2653_adj_1185), .Z(n2752_adj_1047)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1802_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1793_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[20]), 
         .D(n2644_adj_1168), .Z(n2743_adj_966)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1793_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2271_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[11]), 
         .D(n3346_adj_1276), .Z(n23_adj_1277)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2271_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1798_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[15]), 
         .D(n2649_adj_1171), .Z(n2748_adj_1040)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1798_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_2_lut (.A(n1610[31]), .B(n1610[29]), .Z(n33572)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 div_9_i1784_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[29]), 
         .D(n2635_adj_1153), .Z(n2734_adj_650)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1784_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX pwm_cnt_1138__i13 (.D(n50[13]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i13.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i12 (.D(n50[12]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i12.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i11 (.D(n50[11]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i11.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i10 (.D(n50[10]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i10.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i9 (.D(n50[9]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i9.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i8 (.D(n50[8]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i8.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i7 (.D(n50[7]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i7.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i6 (.D(n50[6]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i6.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i5 (.D(n50[5]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i5.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i4 (.D(n50[4]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i4.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i3 (.D(n50[3]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i3.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i2 (.D(n50[2]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i2.GSR = "ENABLED";
    FD1S3IX pwm_cnt_1138__i1 (.D(n50[1]), .CK(fastclk_c), .CD(n14116), 
            .Q(pwm_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_131 (.A(n3327), .B(n34842), .C(n3339), .D(n3344), 
         .Z(n34848)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_131.init = 16'hfffe;
    LUT4 i1_4_lut_adj_132 (.A(n3342), .B(n34838), .C(n34816), .D(n3326), 
         .Z(n34846)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_132.init = 16'hfffe;
    CCU2C div_13_add_1311_15 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[29]), 
          .D0(n1843_adj_1189), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[30]), 
          .D1(n1842_adj_1190), .CIN(n30899), .COUT(n30900), .S0(n2006_adj_2182[29]), 
          .S1(n2006_adj_2182[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1311_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1311_15.INJECT1_0 = "NO";
    defparam div_13_add_1311_15.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_133 (.A(n1944), .B(n2006[27]), .C(n38282), 
         .D(n2042_adj_849), .Z(n35692)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_133.init = 16'hffca;
    LUT4 i1_4_lut_adj_134 (.A(n3332), .B(n3336), .C(n3328), .D(n3343), 
         .Z(n34842)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_134.init = 16'hfffe;
    LUT4 div_13_i1252_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[25]), 
         .D(n1847_adj_1192), .Z(n1946_adj_1128)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1252_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1254_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[23]), 
         .D(n1849_adj_1193), .Z(n1948_adj_1132)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1254_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2073_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[8]), 
         .D(n38216), .Z(n3151_adj_1294)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2073_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_135 (.A(n3341), .B(n3330), .C(n3334), .D(n3345), 
         .Z(n34838)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_135.init = 16'hfffe;
    LUT4 rem_10_i2065_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[16]), 
         .D(n3044_adj_1296), .Z(n3143_adj_1297)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2065_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_136 (.A(n34732), .B(n34782), .C(n1650), .D(n28104), 
         .Z(n28562)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_136.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_137 (.A(n1647), .B(n1648), .C(n1649), .Z(n34732)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_137.init = 16'h8080;
    LUT4 i24153_3_lut (.A(n332), .B(n1653), .C(n1654), .Z(n28104)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24153_3_lut.init = 16'hecec;
    LUT4 div_13_i1055_3_lut (.A(n330), .B(n1610[21]), .C(n28558), .Z(n1653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1055_3_lut.init = 16'hcaca;
    LUT4 div_13_i1056_3_lut (.A(n331), .B(n1610[20]), .C(n28558), .Z(n1654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1056_3_lut.init = 16'hcaca;
    LUT4 div_13_i1054_3_lut (.A(n329), .B(n1610[22]), .C(n28558), .Z(n1652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1054_3_lut.init = 16'hcaca;
    LUT4 div_13_i1049_3_lut (.A(n1350), .B(n1610[27]), .C(n28558), .Z(n1647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1049_3_lut.init = 16'hcaca;
    LUT4 div_13_i1050_3_lut (.A(n1351), .B(n1610[26]), .C(n28558), .Z(n1648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1050_3_lut.init = 16'hcaca;
    LUT4 div_13_i1051_3_lut (.A(n1352), .B(n1610[25]), .C(n28558), .Z(n1649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1051_3_lut.init = 16'hcaca;
    LUT4 div_9_i1786_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[27]), 
         .D(n2637_adj_1166), .Z(n2736_adj_663)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1786_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1052_3_lut (.A(n1353), .B(n1610[24]), .C(n28558), .Z(n1650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1052_3_lut.init = 16'hcaca;
    LUT4 div_13_i1048_3_lut (.A(n1448), .B(n1610[28]), .C(n28558), .Z(n1646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1048_3_lut.init = 16'hcaca;
    LUT4 div_13_i2063_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[18]), 
         .D(n3042_adj_1299), .Z(n3141_adj_730)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2063_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1792_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[21]), 
         .D(n2643_adj_1167), .Z(n2742_adj_762)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1792_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1782_3_lut_rep_238_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[31]), 
         .D(n2633), .Z(n38243)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1782_3_lut_rep_238_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1791_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[22]), 
         .D(n2642_adj_1302), .Z(n2741_adj_1036)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1791_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1796_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[17]), 
         .D(n2647_adj_1169), .Z(n2746_adj_1034)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1796_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2251_3_lut_4_lut (.A(n28512), .B(n13602), .C(n3392[31]), 
         .D(n3326_adj_1304), .Z(n63_adj_1305)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2251_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1788_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[25]), 
         .D(n2639_adj_1164), .Z(n2738_adj_1089)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1788_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_54_i27_2_lut (.A(pwm_cnt[13]), .B(duty0[13]), .Z(n36756)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i27_2_lut.init = 16'h9999;
    LUT4 n3397_bdd_4_lut (.A(n3328_adj_1306), .B(n3330_adj_613), .C(n38173), 
         .D(n3338_adj_1307), .Z(n37487)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3397_bdd_4_lut.init = 16'hfffe;
    LUT4 div_9_i1789_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[24]), 
         .D(n2640_adj_1162), .Z(n2739_adj_1035)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1789_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1783_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[30]), 
         .D(n2634_adj_1163), .Z(n2733_adj_1019)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1783_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32208_4_lut (.A(n38362), .B(n36756), .C(n38364), .D(n36720), 
         .Z(n36935)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i32208_4_lut.init = 16'hbfbb;
    LUT4 div_9_i1799_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[14]), 
         .D(n2650_adj_1173), .Z(n2749_adj_1041)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1799_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1804_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[9]), 
         .D(n342_adj_1184), .Z(n2754_adj_1038)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1804_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_138 (.A(n36286), .B(n2437_adj_1310), .C(n36270), 
         .D(n2445_adj_1311), .Z(n13554)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_138.init = 16'hfffe;
    LUT4 i1_4_lut_adj_139 (.A(n2438_adj_1312), .B(n36282), .C(n36268), 
         .D(n2446_adj_1313), .Z(n36286)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_139.init = 16'hfffe;
    LUT4 div_9_i1803_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[10]), 
         .D(n2654_adj_1186), .Z(n2753_adj_1043)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1803_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2050_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[31]), 
         .D(n3029_adj_1316), .Z(n3128)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2050_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_140 (.A(n2439_adj_1317), .B(n2436_adj_1318), .C(n2435), 
         .D(n2443_adj_1319), .Z(n36282)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_140.init = 16'hfffe;
    LUT4 i1_4_lut_adj_141 (.A(n2447_adj_1320), .B(n28228), .C(n2448_adj_1321), 
         .D(n2449_adj_1322), .Z(n28319)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_141.init = 16'h8000;
    LUT4 i24276_4_lut (.A(n2451_adj_1323), .B(n2450_adj_1324), .C(n27964), 
         .D(n2452_adj_1325), .Z(n28228)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24276_4_lut.init = 16'heccc;
    LUT4 i24014_3_lut (.A(n340_adj_1326), .B(n2453_adj_1327), .C(n2454_adj_1328), 
         .Z(n27964)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24014_3_lut.init = 16'hecec;
    LUT4 div_9_i1794_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[19]), 
         .D(n38252), .Z(n2744_adj_1032)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1794_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1785_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[28]), 
         .D(n2636_adj_1154), .Z(n2735_adj_998)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1785_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24466_4_lut (.A(n1352), .B(n1350), .C(n1351), .D(n28126), 
         .Z(n28420)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24466_4_lut.init = 16'heccc;
    LUT4 div_9_i1795_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[18]), 
         .D(n2646_adj_1157), .Z(n2745_adj_1033)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1795_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24175_3_lut (.A(n329), .B(n1353), .C(n1354), .Z(n28126)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24175_3_lut.init = 16'hecec;
    LUT4 i4847_2_lut (.A(n38[28]), .B(n3556), .Z(n446)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4847_2_lut.init = 16'h8888;
    LUT4 div_9_i1797_3_lut_4_lut (.A(n28544), .B(n13552), .C(n2699_adj_2181[16]), 
         .D(n2648_adj_1170), .Z(n2747_adj_1039)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24586_2_lut_rep_243 (.A(n28432), .B(n13606), .Z(n38248)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24586_2_lut_rep_243.init = 16'heeee;
    LUT4 rem_10_i1784_3_lut_rep_237_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[29]), 
         .D(n2635_adj_1146), .Z(n38242)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1784_3_lut_rep_237_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1786_3_lut_rep_239_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[27]), 
         .D(n2637_adj_1202), .Z(n38244)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1786_3_lut_rep_239_4_lut.init = 16'hf1e0;
    LUT4 i32127_4_lut_4_lut (.A(n38362), .B(n36756), .C(n14_adj_1332), 
         .D(n4), .Z(n26_adj_1333)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i32127_4_lut_4_lut.init = 16'hf4b0;
    LUT4 rem_10_i1802_3_lut_rep_241_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[11]), 
         .D(n2653_adj_1214), .Z(n38246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1802_3_lut_rep_241_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1797_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[16]), 
         .D(n2648_adj_1335), .Z(n2747_adj_824)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32129_4_lut_4_lut (.A(n38366), .B(n36813), .C(n14_adj_1336), 
         .D(n4_adj_1337), .Z(n26_adj_1338)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i32129_4_lut_4_lut.init = 16'hf4b0;
    LUT4 rem_10_i1798_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[15]), 
         .D(n2649_adj_1340), .Z(n2748_adj_911)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1798_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32131_4_lut_4_lut (.A(n38370), .B(n36870), .C(n14_adj_1341), 
         .D(n4_adj_1342), .Z(n26_adj_1178)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32131_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i32133_4_lut_4_lut (.A(n38374), .B(n36927), .C(n14_adj_1343), 
         .D(n4_adj_1344), .Z(n26_adj_842)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32133_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i32135_4_lut_4_lut (.A(n38380), .B(n36747), .C(n20_adj_1345), 
         .D(n6_adj_1346), .Z(n22_adj_653)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i32135_4_lut_4_lut.init = 16'hf4b0;
    LUT4 rem_10_i1782_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[31]), 
         .D(n2633_adj_1348), .Z(n2732_adj_648)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1782_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32200_4_lut_4_lut (.A(n38380), .B(n36743), .C(n36756), .D(n38362), 
         .Z(n36760)) /* synthesis lut_function=(A ((D)+!C)+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i32200_4_lut_4_lut.init = 16'hff4f;
    LUT4 i32137_4_lut_4_lut (.A(n38386), .B(n36804), .C(n20_adj_1349), 
         .D(n6_adj_1350), .Z(n22_adj_626)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i32137_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i32176_4_lut_4_lut (.A(n38386), .B(n36800), .C(n36813), .D(n38366), 
         .Z(n36817)) /* synthesis lut_function=(A ((D)+!C)+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i32176_4_lut_4_lut.init = 16'hff4f;
    LUT4 i32139_4_lut_4_lut (.A(n38392), .B(n36861), .C(n20_adj_1351), 
         .D(n6_adj_1352), .Z(n22_adj_608)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32139_4_lut_4_lut.init = 16'hf4b0;
    LUT4 div_13_i2064_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[17]), 
         .D(n3043_adj_1354), .Z(n3142_adj_684)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2064_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1847_15 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[21]), 
          .D0(n2643_adj_1167), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[22]), 
          .D1(n2642_adj_1302), .CIN(n30740), .COUT(n30741), .S0(n2798_adj_2166[21]), 
          .S1(n2798_adj_2166[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_15.INJECT1_0 = "NO";
    defparam div_9_add_1847_15.INJECT1_1 = "NO";
    LUT4 rem_10_i1799_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[14]), 
         .D(n2650_adj_1356), .Z(n2749_adj_941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1799_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32218_4_lut_4_lut (.A(n38392), .B(n36857), .C(n36870), .D(n38370), 
         .Z(n36874)) /* synthesis lut_function=(A ((D)+!C)+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32218_4_lut_4_lut.init = 16'hff4f;
    LUT4 div_13_i2060_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[21]), 
         .D(n3039_adj_1358), .Z(n3138_adj_661)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2060_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1244_3 (.A0(n38307), .B0(n1808_adj_2179[18]), .C0(n35[18]), 
          .D0(n38293), .A1(n13653), .B1(n28287), .C1(n1808_adj_2179[19]), 
          .D1(n1754_adj_1076), .CIN(n30638), .COUT(n30639), .S0(n1907_adj_2173[18]), 
          .S1(n1907_adj_2173[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_3.INIT0 = 16'hcca0;
    defparam div_9_add_1244_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1244_3.INJECT1_0 = "NO";
    defparam div_9_add_1244_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1804_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[9]), 
         .D(n591), .Z(n2754_adj_945)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1804_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1794_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[19]), 
         .D(n2645_adj_1363), .Z(n2744_adj_822)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1794_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1801_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[12]), 
         .D(n2652_adj_1365), .Z(n2751_adj_950)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1801_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1791_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[22]), 
         .D(n2642_adj_1367), .Z(n2741_adj_780)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1791_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1800_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[13]), 
         .D(n2651_adj_1369), .Z(n2750_adj_943)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1800_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1790_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[23]), 
         .D(n2641_adj_1371), .Z(n2740)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1790_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2073_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[8]), 
         .D(n3052_adj_1373), .Z(n3151)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2073_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32141_4_lut_4_lut (.A(n38398), .B(n36918), .C(n20_adj_1374), 
         .D(n6_adj_1375), .Z(n22)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32141_4_lut_4_lut.init = 16'hf4b0;
    LUT4 rem_10_i1783_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[30]), 
         .D(n2634_adj_1377), .Z(n2733_adj_884)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1783_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32213_4_lut_4_lut (.A(n38398), .B(n36914), .C(n36927), .D(n38374), 
         .Z(n36931)) /* synthesis lut_function=(A ((D)+!C)+!A (B+((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32213_4_lut_4_lut.init = 16'hff4f;
    CCU2C div_9_add_1244_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n39), .D1(n35[17]), 
          .COUT(n30638), .S1(n1907_adj_2173[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1244_1.INIT0 = 16'h0000;
    defparam div_9_add_1244_1.INIT1 = 16'habef;
    defparam div_9_add_1244_1.INJECT1_0 = "NO";
    defparam div_9_add_1244_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1311_13 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[27]), 
          .D0(n1845_adj_1379), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[28]), 
          .D1(n1844_adj_1188), .CIN(n30898), .COUT(n30899), .S0(n2006_adj_2182[27]), 
          .S1(n2006_adj_2182[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1311_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1311_13.INJECT1_0 = "NO";
    defparam div_13_add_1311_13.INJECT1_1 = "NO";
    LUT4 div_13_i2072_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[9]), 
         .D(n3051_adj_1382), .Z(n3150_adj_697)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2072_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1847_13 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[19]), 
          .D0(n38252), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[20]), 
          .D1(n2644_adj_1168), .CIN(n30739), .COUT(n30740), .S0(n2798_adj_2166[19]), 
          .S1(n2798_adj_2166[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_13.INJECT1_0 = "NO";
    defparam div_9_add_1847_13.INJECT1_1 = "NO";
    CCU2C div_9_add_1847_11 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[17]), 
          .D0(n2647_adj_1169), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[18]), 
          .D1(n2646_adj_1157), .CIN(n30738), .COUT(n30739), .S0(n2798_adj_2166[17]), 
          .S1(n2798_adj_2166[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_11.INJECT1_0 = "NO";
    defparam div_9_add_1847_11.INJECT1_1 = "NO";
    CCU2C div_13_add_1311_11 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[25]), 
          .D0(n1847_adj_1192), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[26]), 
          .D1(n1846_adj_1384), .CIN(n30897), .COUT(n30898), .S0(n2006_adj_2182[25]), 
          .S1(n2006_adj_2182[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1311_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1311_11.INJECT1_0 = "NO";
    defparam div_13_add_1311_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1177_15 (.A0(n38305), .B0(GND_net), .C0(n1709_adj_2160[31]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30637), .S0(n1808_adj_2179[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1177_15.INIT1 = 16'h0000;
    defparam div_9_add_1177_15.INJECT1_0 = "NO";
    defparam div_9_add_1177_15.INJECT1_1 = "NO";
    LUT4 div_13_i2065_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[16]), 
         .D(n3044_adj_1386), .Z(n3143)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2065_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1788_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[25]), 
         .D(n2639_adj_1388), .Z(n2738_adj_760)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1788_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1177_13 (.A0(n38305), .B0(GND_net), .C0(n1709_adj_2160[29]), 
          .D0(GND_net), .A1(n38305), .B1(GND_net), .C1(n1709_adj_2160[30]), 
          .D1(GND_net), .CIN(n30636), .COUT(n30637), .S0(n1808_adj_2179[29]), 
          .S1(n1808_adj_2179[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1177_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1177_13.INJECT1_0 = "NO";
    defparam div_9_add_1177_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1311_9 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[23]), 
          .D0(n1849_adj_1193), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[24]), 
          .D1(n1848_adj_1191), .CIN(n30896), .COUT(n30897), .S0(n2006_adj_2182[23]), 
          .S1(n2006_adj_2182[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1311_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1311_9.INJECT1_0 = "NO";
    defparam div_13_add_1311_9.INJECT1_1 = "NO";
    LUT4 rem_10_i1795_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[18]), 
         .D(n2646_adj_1391), .Z(n2745)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1795_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1311_7 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[21]), 
          .D0(n1851_adj_1194), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[22]), 
          .D1(n1850_adj_1195), .CIN(n30895), .COUT(n30896), .S0(n2006_adj_2182[21]), 
          .S1(n2006_adj_2182[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1311_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1311_7.INJECT1_0 = "NO";
    defparam div_13_add_1311_7.INJECT1_1 = "NO";
    LUT4 div_13_i2055_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[26]), 
         .D(n38203), .Z(n3133)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2055_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1311_5 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[19]), 
          .D0(n1853_adj_1200), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[20]), 
          .D1(n1852_adj_1196), .CIN(n30894), .COUT(n30895), .S0(n2006_adj_2182[19]), 
          .S1(n2006_adj_2182[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1311_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1311_5.INJECT1_0 = "NO";
    defparam div_13_add_1311_5.INJECT1_1 = "NO";
    LUT4 div_13_i2068_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[13]), 
         .D(n3047_adj_1398), .Z(n3146_adj_768)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2068_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1796_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[17]), 
         .D(n2647_adj_1400), .Z(n2746_adj_818)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1796_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1847_9 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[15]), 
          .D0(n2649_adj_1171), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[16]), 
          .D1(n2648_adj_1170), .CIN(n30737), .COUT(n30738), .S0(n2798_adj_2166[15]), 
          .S1(n2798_adj_2166[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1847_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1847_9.INJECT1_0 = "NO";
    defparam div_9_add_1847_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1311_3 (.A0(n38283), .B0(n28377), .C0(n1907_adj_2183[17]), 
          .D0(n334_adj_1199), .A1(n38283), .B1(n28377), .C1(n1907_adj_2183[18]), 
          .D1(n1854_adj_1201), .CIN(n30893), .COUT(n30894), .S0(n2006_adj_2182[17]), 
          .S1(n2006_adj_2182[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1311_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1311_3.INJECT1_0 = "NO";
    defparam div_13_add_1311_3.INJECT1_1 = "NO";
    CCU2C div_9_add_1177_11 (.A0(n38305), .B0(GND_net), .C0(n1709_adj_2160[27]), 
          .D0(GND_net), .A1(n38305), .B1(GND_net), .C1(n1709_adj_2160[28]), 
          .D1(n38305), .CIN(n30635), .COUT(n30636), .S0(n1808_adj_2179[27]), 
          .S1(n1808_adj_2179[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1177_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1177_11.INJECT1_0 = "NO";
    defparam div_9_add_1177_11.INJECT1_1 = "NO";
    LUT4 div_13_i2069_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[12]), 
         .D(n3048_adj_1404), .Z(n3147_adj_770)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2069_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2062_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[19]), 
         .D(n38208), .Z(n3140_adj_772)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2062_3_lut_4_lut.init = 16'hf1e0;
    PFUMX pwm_cnt_14__I_0_53_i28 (.BLUT(n12_adj_1406), .ALUT(n26_adj_1338), 
          .C0(n36939), .Z(n28_adj_1407)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    CCU2C div_9_add_1847_7 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[13]), 
          .D0(n2651_adj_1172), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[14]), 
          .D1(n2650_adj_1173), .CIN(n30736), .COUT(n30737), .S0(n2798_adj_2166[13]), 
          .S1(n2798_adj_2166[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1847_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1847_7.INJECT1_0 = "NO";
    defparam div_9_add_1847_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1177_9 (.A0(n38305), .B0(GND_net), .C0(n1709_adj_2160[25]), 
          .D0(n38305), .A1(n38305), .B1(GND_net), .C1(n1709_adj_2160[26]), 
          .D1(GND_net), .CIN(n30634), .COUT(n30635), .S0(n1808_adj_2179[25]), 
          .S1(n1808_adj_2179[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1177_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1177_9.INJECT1_0 = "NO";
    defparam div_9_add_1177_9.INJECT1_1 = "NO";
    CCU2C div_9_add_1847_5 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[11]), 
          .D0(n2653_adj_1185), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[12]), 
          .D1(n2652_adj_1174), .CIN(n30735), .COUT(n30736), .S0(n2798_adj_2166[11]), 
          .S1(n2798_adj_2166[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1847_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1847_5.INJECT1_0 = "NO";
    defparam div_9_add_1847_5.INJECT1_1 = "NO";
    CCU2C div_9_add_1177_7 (.A0(n38305), .B0(GND_net), .C0(n1709_adj_2160[23]), 
          .D0(GND_net), .A1(n38305), .B1(GND_net), .C1(n1709_adj_2160[24]), 
          .D1(GND_net), .CIN(n30633), .COUT(n30634), .S0(n1808_adj_2179[23]), 
          .S1(n1808_adj_2179[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1177_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1177_7.INJECT1_0 = "NO";
    defparam div_9_add_1177_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1311_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n335_adj_1150), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30893), .S1(n2006_adj_2182[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1311_1.INIT0 = 16'h0000;
    defparam div_13_add_1311_1.INIT1 = 16'h555a;
    defparam div_13_add_1311_1.INJECT1_0 = "NO";
    defparam div_13_add_1311_1.INJECT1_1 = "NO";
    LUT4 rem_10_i1785_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[28]), 
         .D(n38250), .Z(n2735_adj_814)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1785_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1803_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[10]), 
         .D(n2654_adj_1413), .Z(n2753_adj_774)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1803_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2414_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3556), 
         .D(n4990[4]), .Z(n197[4])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2414_3_lut_4_lut.init = 16'hfe0e;
    LUT4 rem_10_i1793_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[20]), 
         .D(n2644_adj_1415), .Z(n2743_adj_890)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1793_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_2_lut_rep_347 (.A(distance[10]), .B(distance[13]), .Z(n38352)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_rep_347.init = 16'heeee;
    LUT4 div_13_i2053_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[28]), 
         .D(n3032_adj_1417), .Z(n3131)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2053_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1792_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[21]), 
         .D(n2643_adj_1419), .Z(n2742_adj_892)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1792_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1244_15 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[30]), 
          .D0(n1743_adj_1421), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[31]), 
          .D1(n1742_adj_1423), .CIN(n30891), .S0(n1907_adj_2183[30]), 
          .S1(n1907_adj_2183[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1244_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1244_15.INJECT1_0 = "NO";
    defparam div_13_add_1244_15.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_173 (.A(n3452), .B(n3453), .C(n3451), .Z(n38178)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_3_lut_rep_173.init = 16'h8080;
    CCU2C div_13_add_1244_13 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[28]), 
          .D0(n1745_adj_1425), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[29]), 
          .D1(n38286), .CIN(n30890), .COUT(n30891), .S0(n1907_adj_2183[28]), 
          .S1(n1907_adj_2183[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1244_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1244_13.INJECT1_0 = "NO";
    defparam div_13_add_1244_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1787_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[26]), 
         .D(n2638_adj_1428), .Z(n2737_adj_798)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1787_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32163_2_lut_4_lut (.A(n1), .B(n13790), .C(n89[0]), .D(n12416), 
         .Z(n12429)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i32163_2_lut_4_lut.init = 16'hffdf;
    LUT4 i3_2_lut_rep_348 (.A(distance[14]), .B(distance[12]), .Z(n38353)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut_rep_348.init = 16'heeee;
    CCU2C div_9_add_1177_5 (.A0(n38305), .B0(GND_net), .C0(n1709_adj_2160[21]), 
          .D0(n38305), .A1(n38305), .B1(GND_net), .C1(n1709_adj_2160[22]), 
          .D1(n38305), .CIN(n30632), .COUT(n30633), .S0(n1808_adj_2179[21]), 
          .S1(n1808_adj_2179[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1177_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1177_5.INJECT1_0 = "NO";
    defparam div_9_add_1177_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut (.A(distance[14]), .B(distance[12]), .C(distance[13]), 
         .D(distance[10]), .Z(n34948)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    CCU2C div_13_add_1244_11 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[26]), 
          .D0(n1747_adj_1430), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[27]), 
          .D1(n1746_adj_1432), .CIN(n30889), .COUT(n30890), .S0(n1907_adj_2183[26]), 
          .S1(n1907_adj_2183[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1244_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1244_11.INJECT1_0 = "NO";
    defparam div_13_add_1244_11.INJECT1_1 = "NO";
    LUT4 rem_10_i1789_3_lut_4_lut (.A(n28432), .B(n13606), .C(n2699_adj_2180[24]), 
         .D(n2640_adj_1434), .Z(n2739_adj_816)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1789_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24506_2_lut_rep_244 (.A(n28456), .B(n13625), .Z(n38249)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24506_2_lut_rep_244.init = 16'heeee;
    CCU2C div_13_add_1244_9 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[24]), 
          .D0(n1749_adj_1436), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[25]), 
          .D1(n1748_adj_1438), .CIN(n30888), .COUT(n30889), .S0(n1907_adj_2183[24]), 
          .S1(n1907_adj_2183[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1244_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1244_9.INJECT1_0 = "NO";
    defparam div_13_add_1244_9.INJECT1_1 = "NO";
    CCU2C div_9_add_1847_3 (.A0(n13552), .B0(n28544), .C0(n2699_adj_2181[9]), 
          .D0(n342_adj_1184), .A1(n13552), .B1(n28544), .C1(n2699_adj_2181[10]), 
          .D1(n2654_adj_1186), .CIN(n30734), .COUT(n30735), .S0(n2798_adj_2166[9]), 
          .S1(n2798_adj_2166[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1847_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1847_3.INJECT1_0 = "NO";
    defparam div_9_add_1847_3.INJECT1_1 = "NO";
    LUT4 div_13_i1730_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[16]), 
         .D(n2549), .Z(n2648)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1730_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1177_3 (.A0(n38307), .B0(n1709_adj_2160[19]), .C0(n35[19]), 
          .D0(n38305), .A1(n38305), .B1(GND_net), .C1(n1709_adj_2160[20]), 
          .D1(n38305), .CIN(n30631), .COUT(n30632), .S0(n1808_adj_2179[19]), 
          .S1(n1808_adj_2179[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_3.INIT0 = 16'hcca0;
    defparam div_9_add_1177_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1177_3.INJECT1_0 = "NO";
    defparam div_9_add_1177_3.INJECT1_1 = "NO";
    LUT4 div_13_i1717_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[29]), 
         .D(n2536), .Z(n2635)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1717_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1244_7 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[22]), 
          .D0(n1751_adj_1441), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[23]), 
          .D1(n1750_adj_1443), .CIN(n30887), .COUT(n30888), .S0(n1907_adj_2183[22]), 
          .S1(n1907_adj_2183[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1244_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1244_7.INJECT1_0 = "NO";
    defparam div_13_add_1244_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1177_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n35[18]), 
          .COUT(n30631), .S1(n1808_adj_2179[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1177_1.INIT0 = 16'h0000;
    defparam div_9_add_1177_1.INIT1 = 16'hdfff;
    defparam div_9_add_1177_1.INJECT1_0 = "NO";
    defparam div_9_add_1177_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1847_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n66_adj_9), .D1(n35[8]), 
          .COUT(n30734), .S1(n2798_adj_2166[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1847_1.INIT0 = 16'h0000;
    defparam div_9_add_1847_1.INIT1 = 16'habef;
    defparam div_9_add_1847_1.INJECT1_0 = "NO";
    defparam div_9_add_1847_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1244_5 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[20]), 
          .D0(n1753_adj_724), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[21]), 
          .D1(n38287), .CIN(n30886), .COUT(n30887), .S0(n1907_adj_2183[20]), 
          .S1(n1907_adj_2183[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1244_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1244_5.INJECT1_0 = "NO";
    defparam div_13_add_1244_5.INJECT1_1 = "NO";
    CCU2C div_9_add_1780_23 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[30]), 
          .D0(n2535_adj_1246), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[31]), 
          .D1(n2534_adj_1248), .CIN(n30732), .S0(n2699_adj_2181[30]), 
          .S1(n2699_adj_2181[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_23.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_23.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_23.INJECT1_0 = "NO";
    defparam div_9_add_1780_23.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i4_4_lut_4_lut (.A(pwm_cnt[0]), .B(pwm_cnt[1]), 
         .C(duty1[1]), .D(duty1[0]), .Z(n4_adj_1337)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_14__I_0_53_i4_4_lut_4_lut.init = 16'h7130;
    LUT4 pwm_cnt_14__I_0_52_i4_4_lut_4_lut (.A(pwm_cnt[0]), .B(pwm_cnt[1]), 
         .C(duty2[1]), .D(duty2[0]), .Z(n4_adj_1342)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_14__I_0_52_i4_4_lut_4_lut.init = 16'h7130;
    LUT4 div_13_i2067_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[14]), 
         .D(n3046_adj_1449), .Z(n3145_adj_806)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2067_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1728_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[18]), 
         .D(n2547), .Z(n2646)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1728_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1110_13 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2187[30]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2187[31]), 
          .D1(GND_net), .CIN(n30629), .S0(n1709_adj_2160[30]), .S1(n1709_adj_2160[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_13.INIT0 = 16'h0f1f;
    defparam div_9_add_1110_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1110_13.INJECT1_0 = "NO";
    defparam div_9_add_1110_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1244_3 (.A0(n13638), .B0(n28566), .C0(n1808_adj_2185[18]), 
          .D0(n333_adj_1452), .A1(n13638), .B1(n28566), .C1(n1808_adj_2185[19]), 
          .D1(n1754_adj_1454), .CIN(n30885), .COUT(n30886), .S0(n1907_adj_2183[18]), 
          .S1(n1907_adj_2183[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1244_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1244_3.INJECT1_0 = "NO";
    defparam div_13_add_1244_3.INJECT1_1 = "NO";
    LUT4 div_13_i1729_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[17]), 
         .D(n2548), .Z(n2647)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1729_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1780_21 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[28]), 
          .D0(n2537_adj_1236), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[29]), 
          .D1(n2536_adj_1237), .CIN(n30731), .COUT(n30732), .S0(n2699_adj_2181[28]), 
          .S1(n2699_adj_2181[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_21.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_21.INJECT1_0 = "NO";
    defparam div_9_add_1780_21.INJECT1_1 = "NO";
    CCU2C div_13_add_1244_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n334_adj_1199), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30885), .S1(n1907_adj_2183[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1244_1.INIT0 = 16'h0000;
    defparam div_13_add_1244_1.INIT1 = 16'h555a;
    defparam div_13_add_1244_1.INJECT1_0 = "NO";
    defparam div_13_add_1244_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1177_15 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[31]), 
          .D0(n1643), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30884), .S0(n1808_adj_2185[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1177_15.INIT1 = 16'h0000;
    defparam div_13_add_1177_15.INJECT1_0 = "NO";
    defparam div_13_add_1177_15.INJECT1_1 = "NO";
    CCU2C div_9_add_1780_19 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[26]), 
          .D0(n2539_adj_1235), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[27]), 
          .D1(n2538_adj_1245), .CIN(n30730), .COUT(n30731), .S0(n2699_adj_2181[26]), 
          .S1(n2699_adj_2181[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_19.INJECT1_0 = "NO";
    defparam div_9_add_1780_19.INJECT1_1 = "NO";
    CCU2C div_13_add_1177_13 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[29]), 
          .D0(n1645), .A1(n13640), .B1(n28562), .C1(n1709_adj_2169[30]), 
          .D1(n38294), .CIN(n30883), .COUT(n30884), .S0(n1808_adj_2185[29]), 
          .S1(n1808_adj_2185[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1177_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1177_13.INJECT1_0 = "NO";
    defparam div_13_add_1177_13.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i4_4_lut_4_lut (.A(pwm_cnt[0]), .B(pwm_cnt[1]), 
         .C(duty0[1]), .D(duty0[0]), .Z(n4)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_14__I_0_54_i4_4_lut_4_lut.init = 16'h7130;
    LUT4 div_13_i1725_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[21]), 
         .D(n2544), .Z(n2643)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1725_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1177_11 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[27]), 
          .D0(n1647), .A1(n13640), .B1(n28562), .C1(n1709_adj_2169[28]), 
          .D1(n1646), .CIN(n30882), .COUT(n30883), .S0(n1808_adj_2185[27]), 
          .S1(n1808_adj_2185[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1177_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1177_11.INJECT1_0 = "NO";
    defparam div_13_add_1177_11.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_51_i4_4_lut_4_lut (.A(pwm_cnt[0]), .B(pwm_cnt[1]), 
         .C(duty3[1]), .D(duty3[0]), .Z(n4_adj_1344)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))+!B (C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_14__I_0_51_i4_4_lut_4_lut.init = 16'h7130;
    CCU2C div_13_add_1177_9 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[25]), 
          .D0(n1649), .A1(n13640), .B1(n28562), .C1(n1709_adj_2169[26]), 
          .D1(n1648), .CIN(n30881), .COUT(n30882), .S0(n1808_adj_2185[25]), 
          .S1(n1808_adj_2185[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1177_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1177_9.INJECT1_0 = "NO";
    defparam div_13_add_1177_9.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i7_2_lut_rep_349 (.A(pwm_cnt[3]), .B(duty0[3]), 
         .Z(n38354)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i7_2_lut_rep_349.init = 16'h6666;
    CCU2C div_9_add_1110_11 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2187[28]), 
          .D0(n38305), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2187[29]), 
          .D1(GND_net), .CIN(n30628), .COUT(n30629), .S0(n1709_adj_2160[28]), 
          .S1(n1709_adj_2160[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1110_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1110_11.INJECT1_0 = "NO";
    defparam div_9_add_1110_11.INJECT1_1 = "NO";
    LUT4 i26377_2_lut_rep_170_4_lut (.A(n3452), .B(n3453), .C(n3451), 
         .D(n3450), .Z(n38175)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i26377_2_lut_rep_170_4_lut.init = 16'hff80;
    LUT4 div_13_i2056_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[25]), 
         .D(n3035_adj_1469), .Z(n3134_adj_794)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2056_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_54_i6_3_lut_3_lut (.A(pwm_cnt[3]), .B(duty0[3]), 
         .C(duty0[2]), .Z(n6_adj_1346)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i6_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_13_add_1177_7 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[23]), 
          .D0(n38296), .A1(n13640), .B1(n28562), .C1(n1709_adj_2169[24]), 
          .D1(n1650), .CIN(n30880), .COUT(n30881), .S0(n1808_adj_2185[23]), 
          .S1(n1808_adj_2185[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1177_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1177_7.INJECT1_0 = "NO";
    defparam div_13_add_1177_7.INJECT1_1 = "NO";
    LUT4 div_13_i1716_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[30]), 
         .D(n2535), .Z(n2634)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1716_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1177_5 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[21]), 
          .D0(n1653), .A1(n13640), .B1(n28562), .C1(n1709_adj_2169[22]), 
          .D1(n1652), .CIN(n30879), .COUT(n30880), .S0(n1808_adj_2185[21]), 
          .S1(n1808_adj_2185[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1177_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1177_5.INJECT1_0 = "NO";
    defparam div_13_add_1177_5.INJECT1_1 = "NO";
    LUT4 div_13_i1731_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[15]), 
         .D(n2550), .Z(n2649)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1731_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1722_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[24]), 
         .D(n2541), .Z(n2640)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1722_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2058_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[23]), 
         .D(n3037_adj_1475), .Z(n3136_adj_791)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2058_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1177_3 (.A0(n13640), .B0(n28562), .C0(n1709_adj_2169[19]), 
          .D0(n332), .A1(n13640), .B1(n28562), .C1(n1709_adj_2169[20]), 
          .D1(n1654), .CIN(n30878), .COUT(n30879), .S0(n1808_adj_2185[19]), 
          .S1(n1808_adj_2185[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1177_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1177_3.INJECT1_0 = "NO";
    defparam div_13_add_1177_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1177_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n333_adj_1452), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30878), .S1(n1808_adj_2185[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1177_1.INIT0 = 16'h0000;
    defparam div_13_add_1177_1.INIT1 = 16'h555a;
    defparam div_13_add_1177_1.INJECT1_0 = "NO";
    defparam div_13_add_1177_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1780_17 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[24]), 
          .D0(n2541_adj_1240), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[25]), 
          .D1(n2540_adj_1238), .CIN(n30729), .COUT(n30730), .S0(n2699_adj_2181[24]), 
          .S1(n2699_adj_2181[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_17.INJECT1_0 = "NO";
    defparam div_9_add_1780_17.INJECT1_1 = "NO";
    CCU2C div_13_add_1110_13 (.A0(GND_net), .B0(n28558), .C0(n1610[30]), 
          .D0(GND_net), .A1(GND_net), .B1(n28558), .C1(n1610[31]), .D1(GND_net), 
          .CIN(n30876), .S0(n1709_adj_2169[30]), .S1(n1709_adj_2169[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_13.INIT0 = 16'h0f1f;
    defparam div_13_add_1110_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1110_13.INJECT1_0 = "NO";
    defparam div_13_add_1110_13.INJECT1_1 = "NO";
    CCU2C div_9_add_1780_15 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[22]), 
          .D0(n2543_adj_1247), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[23]), 
          .D1(n2542_adj_1241), .CIN(n30728), .COUT(n30729), .S0(n2699_adj_2181[22]), 
          .S1(n2699_adj_2181[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_15.INJECT1_0 = "NO";
    defparam div_9_add_1780_15.INJECT1_1 = "NO";
    LUT4 div_13_i1733_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[13]), 
         .D(n2552), .Z(n2651)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1733_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1110_11 (.A0(GND_net), .B0(n28558), .C0(n1610[28]), 
          .D0(n1448), .A1(GND_net), .B1(n28558), .C1(n1610[29]), .D1(GND_net), 
          .CIN(n30875), .COUT(n30876), .S0(n1709_adj_2169[28]), .S1(n1709_adj_2169[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1110_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1110_11.INJECT1_0 = "NO";
    defparam div_13_add_1110_11.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i7_2_lut_rep_350 (.A(pwm_cnt[3]), .B(duty1[3]), 
         .Z(n38355)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i7_2_lut_rep_350.init = 16'h6666;
    LUT4 div_13_i1736_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[10]), 
         .D(n341_adj_605), .Z(n2654)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1736_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2070_3_lut_4_lut (.A(n28518), .B(n13617), .C(n3095_adj_2176[11]), 
         .D(n3049_adj_1483), .Z(n3148_adj_810)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2070_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_53_i6_3_lut_3_lut (.A(pwm_cnt[3]), .B(duty1[3]), 
         .C(duty1[2]), .Z(n6_adj_1350)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i6_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1780_13 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[20]), 
          .D0(n2545_adj_1233), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[21]), 
          .D1(n2544_adj_1239), .CIN(n30727), .COUT(n30728), .S0(n2699_adj_2181[20]), 
          .S1(n2699_adj_2181[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_13.INJECT1_0 = "NO";
    defparam div_9_add_1780_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1110_9 (.A0(GND_net), .B0(n28558), .C0(n1610[26]), 
          .D0(n1351), .A1(GND_net), .B1(n28558), .C1(n1610[27]), .D1(n1350), 
          .CIN(n30874), .COUT(n30875), .S0(n1709_adj_2169[26]), .S1(n1709_adj_2169[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1110_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1110_9.INJECT1_0 = "NO";
    defparam div_13_add_1110_9.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_142 (.A(n14790), .B(n197[14]), .C(n89[0]), .Z(duty2_14__N_473[14])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i1_3_lut_adj_142.init = 16'ha8a8;
    LUT4 div_13_i1724_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[22]), 
         .D(n2543), .Z(n2642)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1724_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1110_7 (.A0(GND_net), .B0(n28558), .C0(n1610[24]), 
          .D0(n1353), .A1(GND_net), .B1(n28558), .C1(n1610[25]), .D1(n1352), 
          .CIN(n30873), .COUT(n30874), .S0(n1709_adj_2169[24]), .S1(n1709_adj_2169[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1110_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1110_7.INJECT1_0 = "NO";
    defparam div_13_add_1110_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1110_5 (.A0(GND_net), .B0(n28558), .C0(n1610[22]), 
          .D0(n329), .A1(GND_net), .B1(n28558), .C1(n1610[23]), .D1(n1354), 
          .CIN(n30872), .COUT(n30873), .S0(n1709_adj_2169[22]), .S1(n1709_adj_2169[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1110_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1110_5.INJECT1_0 = "NO";
    defparam div_13_add_1110_5.INJECT1_1 = "NO";
    CCU2C div_9_add_1780_11 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[18]), 
          .D0(n2547_adj_1249), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[19]), 
          .D1(n2546_adj_1234), .CIN(n30726), .COUT(n30727), .S0(n2699_adj_2181[18]), 
          .S1(n2699_adj_2181[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_11.INJECT1_0 = "NO";
    defparam div_9_add_1780_11.INJECT1_1 = "NO";
    LUT4 div_13_i1715_3_lut_rep_236_4_lut (.A(n28456), .B(n13625), .C(n2600[31]), 
         .D(n2534), .Z(n38241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1715_3_lut_rep_236_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1734_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[12]), 
         .D(n2553), .Z(n2652)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1734_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i77_3_lut (.A(n14790), .B(n197[13]), .C(n89[0]), .Z(duty2_14__N_473[13])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i77_3_lut.init = 16'ha8a8;
    CCU2C div_9_add_1780_9 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[16]), 
          .D0(n2549_adj_1251), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[17]), 
          .D1(n2548_adj_1250), .CIN(n30725), .COUT(n30726), .S0(n2699_adj_2181[16]), 
          .S1(n2699_adj_2181[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1780_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1780_9.INJECT1_0 = "NO";
    defparam div_9_add_1780_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_143 (.A(n38307), .B(n89[0]), .C(n4540[24]), .D(n12416), 
         .Z(n36350)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;
    defparam i1_4_lut_adj_143.init = 16'hffec;
    CCU2C div_13_add_1110_3 (.A0(GND_net), .B0(n28558), .C0(n1610[20]), 
          .D0(n331), .A1(GND_net), .B1(n28558), .C1(n1610[21]), .D1(n330), 
          .CIN(n30871), .COUT(n30872), .S0(n1709_adj_2169[20]), .S1(n1709_adj_2169[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1110_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1110_3.INJECT1_0 = "NO";
    defparam div_13_add_1110_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n332), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30871), .S1(n1709_adj_2169[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1110_1.INIT0 = 16'h0000;
    defparam div_13_add_1110_1.INIT1 = 16'h555a;
    defparam div_13_add_1110_1.INJECT1_0 = "NO";
    defparam div_13_add_1110_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1780_7 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[14]), 
          .D0(n2551_adj_1259), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[15]), 
          .D1(n2550_adj_1260), .CIN(n30724), .COUT(n30725), .S0(n2699_adj_2181[14]), 
          .S1(n2699_adj_2181[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1780_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1780_7.INJECT1_0 = "NO";
    defparam div_9_add_1780_7.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_144 (.A(n14790), .B(n197[8]), .C(n89[0]), .Z(duty2_14__N_473[8])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i1_3_lut_adj_144.init = 16'ha8a8;
    CCU2C div_9_add_1780_5 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[12]), 
          .D0(n2553_adj_1272), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[13]), 
          .D1(n2552_adj_1261), .CIN(n30723), .COUT(n30724), .S0(n2699_adj_2181[12]), 
          .S1(n2699_adj_2181[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1780_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1780_5.INJECT1_0 = "NO";
    defparam div_9_add_1780_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_145 (.A(n14790), .B(n197[7]), .C(n89[0]), .Z(duty2_14__N_473[7])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i1_3_lut_adj_145.init = 16'ha8a8;
    LUT4 div_13_i1727_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[19]), 
         .D(n2546), .Z(n2645)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1727_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_52_i7_2_lut_rep_351 (.A(pwm_cnt[3]), .B(duty2[3]), 
         .Z(n38356)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i7_2_lut_rep_351.init = 16'h6666;
    LUT4 rem_10_i2274_3_lut_rep_174 (.A(n3349), .B(n3392_adj_2163[8]), .C(n3359), 
         .Z(n38179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2274_3_lut_rep_174.init = 16'hcaca;
    LUT4 div_13_i1732_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[14]), 
         .D(n2551), .Z(n2650)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1732_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_52_i6_3_lut_3_lut (.A(pwm_cnt[3]), .B(duty2[3]), 
         .C(duty2[2]), .Z(n6_adj_1352)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_51_i7_2_lut_rep_352 (.A(pwm_cnt[3]), .B(duty3[3]), 
         .Z(n38357)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i7_2_lut_rep_352.init = 16'h6666;
    LUT4 div_13_i1735_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[11]), 
         .D(n2554), .Z(n2653)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1735_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i78_3_lut (.A(n14790), .B(n197[5]), .C(n89[0]), .Z(duty2_14__N_473[5])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i78_3_lut.init = 16'ha8a8;
    LUT4 div_13_i2409_3_lut_4_lut (.A(n28456), .B(n13625), .C(n3556), 
         .D(n4990[9]), .Z(n197[9])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2409_3_lut_4_lut.init = 16'hfe0e;
    LUT4 pwm_cnt_14__I_0_51_i6_3_lut_3_lut (.A(pwm_cnt[3]), .B(duty3[3]), 
         .C(duty3[2]), .Z(n6_adj_1375)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i6_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_3_lut_adj_146 (.A(n14790), .B(n197[2]), .C(n89[0]), .Z(duty2_14__N_473[2])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i1_3_lut_adj_146.init = 16'ha8a8;
    LUT4 i1_3_lut_adj_147 (.A(n14790), .B(n197[1]), .C(n89[0]), .Z(duty2_14__N_473[1])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i1_3_lut_adj_147.init = 16'ha8a8;
    LUT4 i1_2_lut_4_lut_adj_148 (.A(n3152), .B(n3194[7]), .C(n38197), 
         .D(n3252), .Z(n35786)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_148.init = 16'hca00;
    LUT4 select_844_Select_8_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[8]), .Z(duty1_14__N_458[8])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_8_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    LUT4 i24636_2_lut_rep_192 (.A(n28588), .B(n13547), .Z(n38197)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24636_2_lut_rep_192.init = 16'heeee;
    LUT4 div_9_i2141_3_lut_rep_191_4_lut (.A(n28588), .B(n13547), .C(n3194[7]), 
         .D(n3152), .Z(n38196)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2141_3_lut_rep_191_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_0_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[0]), .Z(duty1_14__N_458[0])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_0_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    CCU2C div_13_add_1043_13 (.A0(GND_net), .B0(GND_net), .C0(n1511[31]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30870), .S0(n1610[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_13.INIT0 = 16'h0f1f;
    defparam div_13_add_1043_13.INIT1 = 16'h0000;
    defparam div_13_add_1043_13.INJECT1_0 = "NO";
    defparam div_13_add_1043_13.INJECT1_1 = "NO";
    LUT4 div_13_i1723_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[23]), 
         .D(n2542), .Z(n2641)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1723_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1721_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[25]), 
         .D(n2540), .Z(n2639)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1721_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1719_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[27]), 
         .D(n2538), .Z(n2637)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1719_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1726_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[20]), 
         .D(n2545), .Z(n2644)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1726_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1720_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[26]), 
         .D(n2539), .Z(n2638)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1720_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1718_3_lut_4_lut (.A(n28456), .B(n13625), .C(n2600[28]), 
         .D(n2537), .Z(n2636)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1718_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10126_3_lut_then_4_lut (.A(n38[26]), .B(n3556), .C(n38[28]), 
         .D(n6_adj_1495), .Z(n38408)) /* synthesis lut_function=(!(A (B (C (D)))+!A !((C (D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i10126_3_lut_then_4_lut.init = 16'h7bbb;
    LUT4 i10126_3_lut_else_4_lut (.A(n38[26]), .B(n3556), .C(n38[28]), 
         .D(n6_adj_1495), .Z(n38407)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i10126_3_lut_else_4_lut.init = 16'h4888;
    LUT4 div_9_i2127_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[21]), 
         .D(n3138), .Z(n3237)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2127_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1780_3 (.A0(n13553), .B0(n28331), .C0(n2600_adj_2186[10]), 
          .D0(n341), .A1(n13553), .B1(n28331), .C1(n2600_adj_2186[11]), 
          .D1(n2554_adj_1273), .CIN(n30722), .COUT(n30723), .S0(n2699_adj_2181[10]), 
          .S1(n2699_adj_2181[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1780_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1780_3.INJECT1_0 = "NO";
    defparam div_9_add_1780_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_149 (.A(n2537_adj_1498), .B(n2600_adj_2188[28]), 
         .C(n38251), .D(n2644_adj_1415), .Z(n35636)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_149.init = 16'hffca;
    LUT4 div_13_i1926_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[21]), 
         .D(n2841_adj_616), .Z(n2940_adj_1501)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1926_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1652_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[27]), 
         .D(n2439), .Z(n2538)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1652_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2140_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[8]), 
         .D(n38202), .Z(n3250_adj_554)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2140_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1043_11 (.A0(GND_net), .B0(GND_net), .C0(n1511[29]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1511[30]), 
          .D1(GND_net), .CIN(n30869), .COUT(n30870), .S0(n1610[29]), 
          .S1(n1610[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1043_11.INIT1 = 16'h0f1f;
    defparam div_13_add_1043_11.INJECT1_0 = "NO";
    defparam div_13_add_1043_11.INJECT1_1 = "NO";
    LUT4 div_13_i1258_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[19]), 
         .D(n1853_adj_1200), .Z(n1952_adj_1145)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1258_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_150 (.A(n1745_adj_1502), .B(n1808[28]), .C(n38295), 
         .D(n1841), .Z(n35746)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_150.init = 16'hffca;
    CCU2C div_13_add_1043_9 (.A0(GND_net), .B0(GND_net), .C0(n1511[27]), 
          .D0(n1350), .A1(GND_net), .B1(GND_net), .C1(n1511[28]), .D1(n1448), 
          .CIN(n30868), .COUT(n30869), .S0(n1610[27]), .S1(n1610[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1043_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1043_9.INJECT1_0 = "NO";
    defparam div_13_add_1043_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_151 (.A(n1753), .B(n1808[20]), .C(n38295), 
         .D(n1851), .Z(n34788)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_151.init = 16'hca00;
    LUT4 i1_4_lut_adj_152 (.A(n1709[26]), .B(n5_adj_1503), .C(n1709[25]), 
         .D(n1749), .Z(n28090)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_152.init = 16'h8000;
    CCU2C div_9_add_1780_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[9]), .D1(duty0_14__N_426[7]), 
          .COUT(n30722), .S1(n2699_adj_2181[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1780_1.INIT0 = 16'h0000;
    defparam div_9_add_1780_1.INIT1 = 16'h04bf;
    defparam div_9_add_1780_1.INJECT1_0 = "NO";
    defparam div_9_add_1780_1.INJECT1_1 = "NO";
    LUT4 i24342_2_lut_rep_288 (.A(n28287), .B(n13653), .Z(n38293)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24342_2_lut_rep_288.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_153 (.A(n38259), .B(n4540[10]), .C(n38307), 
         .D(n89[9]), .Z(n35900)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_153.init = 16'hffca;
    LUT4 select_844_Select_7_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[7]), .Z(duty1_14__N_458[7])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_7_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    PFUMX i32292 (.BLUT(n37596), .ALUT(n37595), .C0(n38307), .Z(n37597));
    LUT4 div_13_i1663_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[16]), 
         .D(n2450), .Z(n2549)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1663_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24338_2_lut_rep_163 (.A(n28267), .B(n13608), .Z(n38168)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24338_2_lut_rep_163.init = 16'heeee;
    LUT4 div_13_i1927_3_lut_rep_208_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[20]), 
         .D(n2842_adj_620), .Z(n38213)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1927_3_lut_rep_208_4_lut.init = 16'hf1e0;
    PFUMX pwm_cnt_14__I_0_54_i28 (.BLUT(n12_adj_1506), .ALUT(n26_adj_1333), 
          .C0(n36935), .Z(n28_adj_1507)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    LUT4 div_9_i2137_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[11]), 
         .D(n3148), .Z(n3247)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2137_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_5_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[5]), .Z(duty1_14__N_458[5])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_5_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    LUT4 div_13_i2271_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[11]), 
         .D(n3346_adj_1509), .Z(n23_adj_1510)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2271_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1110_9 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2187[26]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2187[27]), 
          .D1(GND_net), .CIN(n30627), .COUT(n30628), .S0(n1709_adj_2160[26]), 
          .S1(n1709_adj_2160[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1110_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1110_9.INJECT1_0 = "NO";
    defparam div_9_add_1110_9.INJECT1_1 = "NO";
    LUT4 div_13_i1650_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[29]), 
         .D(n2437), .Z(n2536)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1650_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2139_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[9]), 
         .D(n3150), .Z(n3249)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2139_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2119_3_lut_rep_185_4_lut (.A(n28588), .B(n13547), .C(n3194[29]), 
         .D(n3130), .Z(n38190)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2119_3_lut_rep_185_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1661_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[18]), 
         .D(n2448), .Z(n2547)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1661_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1937_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[10]), 
         .D(n2852), .Z(n2951_adj_1514)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1937_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1179_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[31]), 
         .D(n1742), .Z(n1841_adj_874)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1179_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1043_7 (.A0(GND_net), .B0(GND_net), .C0(n1511[25]), 
          .D0(n1352), .A1(GND_net), .B1(GND_net), .C1(n1511[26]), .D1(n1351), 
          .CIN(n30867), .COUT(n30868), .S0(n1610[25]), .S1(n1610[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1043_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1043_7.INJECT1_0 = "NO";
    defparam div_13_add_1043_7.INJECT1_1 = "NO";
    LUT4 div_13_i2267_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[15]), 
         .D(n3342_adj_1516), .Z(n31_adj_1517)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2267_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1662_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[17]), 
         .D(n2449), .Z(n2548)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1662_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_2_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[2]), .Z(duty1_14__N_458[2])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_2_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    CCU2C div_9_add_1110_7 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2187[24]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2187[25]), 
          .D1(n38305), .CIN(n30626), .COUT(n30627), .S0(n1709_adj_2160[24]), 
          .S1(n1709_adj_2160[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1110_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1110_7.INJECT1_0 = "NO";
    defparam div_9_add_1110_7.INJECT1_1 = "NO";
    LUT4 div_13_i2261_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[21]), 
         .D(n3336_adj_1521), .Z(n43_adj_1522)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2261_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1658_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[21]), 
         .D(n2445), .Z(n2544)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1658_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1110_5 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2187[22]), 
          .D0(n38305), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2187[23]), 
          .D1(GND_net), .CIN(n30625), .COUT(n30626), .S0(n1709_adj_2160[22]), 
          .S1(n1709_adj_2160[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1110_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1110_5.INJECT1_0 = "NO";
    defparam div_9_add_1110_5.INJECT1_1 = "NO";
    CCU2C div_13_add_1043_5 (.A0(GND_net), .B0(GND_net), .C0(n1511[23]), 
          .D0(n1354), .A1(GND_net), .B1(GND_net), .C1(n1511[24]), .D1(n1353), 
          .CIN(n30866), .COUT(n30867), .S0(n1610[23]), .S1(n1610[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1043_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1043_5.INJECT1_0 = "NO";
    defparam div_13_add_1043_5.INJECT1_1 = "NO";
    LUT4 div_13_i1657_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[22]), 
         .D(n2444), .Z(n2543)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1657_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2144_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[4]), 
         .D(n347), .Z(n3254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2144_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1043_3 (.A0(GND_net), .B0(GND_net), .C0(n1511[21]), 
          .D0(n330), .A1(GND_net), .B1(GND_net), .C1(n1511[22]), .D1(n329), 
          .CIN(n30865), .COUT(n30866), .S0(n1610[21]), .S1(n1610[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1043_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1043_3.INJECT1_0 = "NO";
    defparam div_13_add_1043_3.INJECT1_1 = "NO";
    LUT4 i10130_3_lut_then_4_lut (.A(n38[24]), .B(n3556), .C(n38[28]), 
         .D(n328), .Z(n38411)) /* synthesis lut_function=(!(A (B (C (D)))+!A !((C (D))+!B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i10130_3_lut_then_4_lut.init = 16'h7bbb;
    LUT4 div_13_i1664_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[15]), 
         .D(n2451), .Z(n2550)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1664_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3359_bdd_4_lut (.A(n38181), .B(n3343_adj_1525), .C(n3337_adj_1526), 
         .D(n3332_adj_1527), .Z(n37665)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3359_bdd_4_lut.init = 16'hfffe;
    LUT4 pwm_cnt_14__I_0_54_i11_2_lut_rep_356 (.A(pwm_cnt[5]), .B(duty0[5]), 
         .Z(n38361)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i11_2_lut_rep_356.init = 16'h6666;
    LUT4 select_842_Select_14_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[14]), 
         .D(n2983), .Z(duty0_14__N_410[14])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_14_i4_3_lut_4_lut.init = 16'hff10;
    CCU2C div_13_add_1043_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n331), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30865), .S1(n1610[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1043_1.INIT0 = 16'h0000;
    defparam div_13_add_1043_1.INIT1 = 16'h555a;
    defparam div_13_add_1043_1.INJECT1_0 = "NO";
    defparam div_13_add_1043_1.INJECT1_1 = "NO";
    LUT4 div_13_i1655_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[24]), 
         .D(n2442), .Z(n2541)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1655_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10130_3_lut_else_4_lut (.A(n38[24]), .B(n3556), .C(n38[28]), 
         .D(n328), .Z(n38410)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i10130_3_lut_else_4_lut.init = 16'h4888;
    LUT4 div_9_i1180_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[30]), 
         .D(n1743), .Z(n1842_adj_957)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2143_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[5]), 
         .D(n3154), .Z(n3253)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2143_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2117_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[31]), 
         .D(n3128_adj_1528), .Z(n3227)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_154 (.A(n3349), .B(n3392_adj_2163[8]), .C(n3359), 
         .D(n3449), .Z(n34936)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_154.init = 16'hca00;
    LUT4 i1_4_lut_adj_155 (.A(n1750), .B(n1709[22]), .C(n7_adj_1529), 
         .D(n1709[21]), .Z(n5_adj_1503)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_155.init = 16'heaaa;
    CCU2C div_9_add_1110_3 (.A0(n38307), .B0(n1610_adj_2187[20]), .C0(n35[19]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2187[21]), 
          .D1(n38305), .CIN(n30624), .COUT(n30625), .S0(n1709_adj_2160[20]), 
          .S1(n1709_adj_2160[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_3.INIT0 = 16'hcca0;
    defparam div_9_add_1110_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1110_3.INJECT1_0 = "NO";
    defparam div_9_add_1110_3.INJECT1_1 = "NO";
    LUT4 select_844_Select_13_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[13]), .Z(duty1_14__N_458[13])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_13_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    CCU2C div_9_add_1713_23 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[31]), 
          .D0(n2435), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30721), .S0(n2600_adj_2186[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_23.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_23.INIT1 = 16'h0000;
    defparam div_9_add_1713_23.INJECT1_0 = "NO";
    defparam div_9_add_1713_23.INJECT1_1 = "NO";
    LUT4 select_844_Select_14_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[14]), .Z(duty1_14__N_458[14])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_14_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    LUT4 pwm_cnt_14__I_0_54_i29_2_lut_rep_357 (.A(pwm_cnt[14]), .B(duty0[14]), 
         .Z(n38362)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i29_2_lut_rep_357.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_54_i14_3_lut_3_lut (.A(pwm_cnt[14]), .B(duty0[14]), 
         .C(duty0[13]), .Z(n14_adj_1332)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i14_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_54_i13_2_lut_rep_358 (.A(pwm_cnt[6]), .B(duty0[6]), 
         .Z(n38363)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i13_2_lut_rep_358.init = 16'h6666;
    CCU2C div_9_add_1110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), 
          .COUT(n30624), .S1(n1709_adj_2160[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1110_1.INIT0 = 16'h0000;
    defparam div_9_add_1110_1.INIT1 = 16'hdfff;
    defparam div_9_add_1110_1.INJECT1_0 = "NO";
    defparam div_9_add_1110_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_156 (.A(n1709[20]), .B(n38306), .C(n1709[19]), .D(n582), 
         .Z(n7_adj_1529)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_156.init = 16'heaaa;
    CCU2C div_9_add_1043_13 (.A0(n38305), .B0(n1412[31]), .C0(n1511_adj_2191[31]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30623), .S0(n1610_adj_2187[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_13.INIT0 = 16'h0fff;
    defparam div_9_add_1043_13.INIT1 = 16'h0000;
    defparam div_9_add_1043_13.INJECT1_0 = "NO";
    defparam div_9_add_1043_13.INJECT1_1 = "NO";
    CCU2C div_9_add_1043_11 (.A0(n38305), .B0(n1412[29]), .C0(n1511_adj_2191[29]), 
          .D0(GND_net), .A1(n38305), .B1(n1412[30]), .C1(n1511_adj_2191[30]), 
          .D1(GND_net), .CIN(n30622), .COUT(n30623), .S0(n1610_adj_2187[29]), 
          .S1(n1610_adj_2187[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_11.INIT0 = 16'h0fff;
    defparam div_9_add_1043_11.INIT1 = 16'h0fff;
    defparam div_9_add_1043_11.INJECT1_0 = "NO";
    defparam div_9_add_1043_11.INJECT1_1 = "NO";
    LUT4 i31884_2_lut_3_lut_4_lut (.A(pwm_cnt[6]), .B(duty0[6]), .C(duty0[5]), 
         .D(pwm_cnt[5]), .Z(n36720)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i31884_2_lut_3_lut_4_lut.init = 16'h9009;
    CCU2C div_13_add_976_11 (.A0(n30262), .B0(n28420), .C0(n446), .D0(n1412_adj_2192[30]), 
          .A1(n30262), .B1(n446), .C1(n28420), .D1(n1412_adj_2192[31]), 
          .CIN(n30863), .S0(n1511[30]), .S1(n1511[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_976_11.INIT0 = 16'hffff;
    defparam div_13_add_976_11.INIT1 = 16'hffff;
    defparam div_13_add_976_11.INJECT1_0 = "NO";
    defparam div_13_add_976_11.INJECT1_1 = "NO";
    CCU2C div_9_add_1713_21 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[29]), 
          .D0(n2437_adj_1310), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[30]), 
          .D1(n2436_adj_1318), .CIN(n30720), .COUT(n30721), .S0(n2600_adj_2186[29]), 
          .S1(n2600_adj_2186[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_21.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_21.INJECT1_0 = "NO";
    defparam div_9_add_1713_21.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i10_3_lut_3_lut (.A(pwm_cnt[6]), .B(duty0[6]), 
         .C(duty0[5]), .Z(n10_adj_1540)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i10_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_54_i15_2_lut_rep_359 (.A(pwm_cnt[7]), .B(duty0[7]), 
         .Z(n38364)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i15_2_lut_rep_359.init = 16'h6666;
    LUT4 div_13_i2256_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[26]), 
         .D(n38172), .Z(n53_adj_1542)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2256_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_54_i12_3_lut_3_lut (.A(pwm_cnt[7]), .B(duty0[7]), 
         .C(n10_adj_1540), .Z(n12_adj_1506)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i12_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1043_9 (.A0(n38305), .B0(n1412[27]), .C0(n1511_adj_2191[27]), 
          .D0(GND_net), .A1(n1412[28]), .B1(n1511_adj_2191[28]), .C1(GND_net), 
          .D1(n38305), .CIN(n30621), .COUT(n30622), .S0(n1610_adj_2187[27]), 
          .S1(n1610_adj_2187[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_9.INIT0 = 16'hf000;
    defparam div_9_add_1043_9.INIT1 = 16'hcfc0;
    defparam div_9_add_1043_9.INJECT1_0 = "NO";
    defparam div_9_add_1043_9.INJECT1_1 = "NO";
    LUT4 div_13_i1667_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[12]), 
         .D(n2454), .Z(n2553)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1667_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1918_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[29]), 
         .D(n38219), .Z(n2932_adj_1546)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1918_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2280_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[2]), 
         .D(n349), .Z(n3454_adj_1548)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2280_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1189_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[21]), 
         .D(n1752_adj_1270), .Z(n1851_adj_963)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1189_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1934_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[13]), 
         .D(n2849_adj_631), .Z(n2948_adj_1550)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1934_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1186_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[24]), 
         .D(n1749_adj_1212), .Z(n1848_adj_959)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1186_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10128_3_lut_then_4_lut (.A(n38[25]), .B(n3556), .C(n38[28]), 
         .D(n30240), .Z(n38414)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(B ((D)+!C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i10128_3_lut_then_4_lut.init = 16'hbb7b;
    LUT4 i10128_3_lut_else_4_lut (.A(n38[25]), .B(n3556), .C(n38[28]), 
         .D(n30240), .Z(n38413)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(((D)+!C)+!B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i10128_3_lut_else_4_lut.init = 16'h8848;
    LUT4 pwm_cnt_14__I_0_53_i11_2_lut_rep_360 (.A(pwm_cnt[5]), .B(duty1[5]), 
         .Z(n38365)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i11_2_lut_rep_360.init = 16'h6666;
    LUT4 div_13_i1935_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[12]), 
         .D(n2850_adj_636), .Z(n2949_adj_1552)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1935_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_53_i29_2_lut_rep_361 (.A(pwm_cnt[14]), .B(duty1[14]), 
         .Z(n38366)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i29_2_lut_rep_361.init = 16'h6666;
    CCU2C div_9_add_1713_19 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[27]), 
          .D0(n2439_adj_1317), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[28]), 
          .D1(n2438_adj_1312), .CIN(n30719), .COUT(n30720), .S0(n2600_adj_2186[27]), 
          .S1(n2600_adj_2186[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_19.INJECT1_0 = "NO";
    defparam div_9_add_1713_19.INJECT1_1 = "NO";
    LUT4 div_9_i1185_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[25]), 
         .D(n38297), .Z(n1847_adj_958)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1920_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[27]), 
         .D(n2835_adj_619), .Z(n2934_adj_1556)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1920_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2278_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[4]), 
         .D(n3353_adj_1558), .Z(n3452_adj_1559)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2278_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2259_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[23]), 
         .D(n3334_adj_1561), .Z(n47)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2259_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_53_i14_3_lut_3_lut (.A(pwm_cnt[14]), .B(duty1[14]), 
         .C(duty1[13]), .Z(n14_adj_1336)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i14_3_lut_3_lut.init = 16'hd4d4;
    FD1S3JX duty3_i14 (.D(duty3_14__N_488[14]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i14.GSR = "DISABLED";
    FD1S3JX duty3_i13 (.D(duty3_14__N_488[13]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i13.GSR = "DISABLED";
    FD1S3IX duty3_i12 (.D(n197[12]), .CK(fastclk_c), .CD(n12429), .Q(duty3[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i12.GSR = "DISABLED";
    FD1S3IX duty3_i11 (.D(n197[11]), .CK(fastclk_c), .CD(n12429), .Q(duty3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i11.GSR = "DISABLED";
    FD1S3IX duty3_i10 (.D(n197[10]), .CK(fastclk_c), .CD(n12429), .Q(duty3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i10.GSR = "DISABLED";
    FD1S3IX duty3_i9 (.D(n197[9]), .CK(fastclk_c), .CD(n12429), .Q(duty3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i9.GSR = "DISABLED";
    FD1S3JX duty3_i8 (.D(duty3_14__N_488[8]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i8.GSR = "DISABLED";
    FD1S3JX duty3_i7 (.D(duty3_14__N_488[7]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i7.GSR = "DISABLED";
    FD1S3IX duty3_i6 (.D(n197[6]), .CK(fastclk_c), .CD(n12429), .Q(duty3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i6.GSR = "DISABLED";
    FD1S3JX duty3_i5 (.D(duty3_14__N_488[5]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i5.GSR = "DISABLED";
    FD1S3IX duty3_i4 (.D(n197[4]), .CK(fastclk_c), .CD(n12429), .Q(duty3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i4.GSR = "DISABLED";
    FD1S3IX duty3_i3 (.D(n197[3]), .CK(fastclk_c), .CD(n12429), .Q(duty3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i3.GSR = "DISABLED";
    FD1S3JX duty3_i2 (.D(duty3_14__N_488[2]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i2.GSR = "DISABLED";
    FD1S3JX duty3_i1 (.D(duty3_14__N_488[1]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty3_i1.GSR = "DISABLED";
    FD1S3JX duty2_i14 (.D(duty2_14__N_473[14]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i14.GSR = "DISABLED";
    FD1S3JX duty2_i13 (.D(duty2_14__N_473[13]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i13.GSR = "DISABLED";
    FD1S3IX duty2_i12 (.D(n197[12]), .CK(fastclk_c), .CD(n13642), .Q(duty2[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i12.GSR = "DISABLED";
    FD1S3IX duty2_i11 (.D(n197[11]), .CK(fastclk_c), .CD(n13642), .Q(duty2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i11.GSR = "DISABLED";
    FD1S3IX duty2_i10 (.D(n197[10]), .CK(fastclk_c), .CD(n13642), .Q(duty2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i10.GSR = "DISABLED";
    FD1S3IX duty2_i9 (.D(n197[9]), .CK(fastclk_c), .CD(n13642), .Q(duty2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i9.GSR = "DISABLED";
    FD1S3JX duty2_i8 (.D(duty2_14__N_473[8]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i8.GSR = "DISABLED";
    FD1S3JX duty2_i7 (.D(duty2_14__N_473[7]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i7.GSR = "DISABLED";
    FD1S3IX duty2_i6 (.D(n197[6]), .CK(fastclk_c), .CD(n13642), .Q(duty2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i6.GSR = "DISABLED";
    FD1S3JX duty2_i5 (.D(duty2_14__N_473[5]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i5.GSR = "DISABLED";
    FD1S3IX duty2_i4 (.D(n197[4]), .CK(fastclk_c), .CD(n13642), .Q(duty2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i4.GSR = "DISABLED";
    FD1S3IX duty2_i3 (.D(n197[3]), .CK(fastclk_c), .CD(n13642), .Q(duty2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i3.GSR = "DISABLED";
    FD1S3JX duty2_i2 (.D(duty2_14__N_473[2]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i2.GSR = "DISABLED";
    FD1S3JX duty2_i1 (.D(duty2_14__N_473[1]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty2_i1.GSR = "DISABLED";
    FD1S3JX duty1_i14 (.D(duty1_14__N_458[14]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i14.GSR = "DISABLED";
    FD1S3JX duty1_i13 (.D(duty1_14__N_458[13]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i13.GSR = "DISABLED";
    FD1S3IX duty1_i12 (.D(duty1_14__N_458[12]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i12.GSR = "DISABLED";
    LUT4 pwm_cnt_14__I_0_53_i13_2_lut_rep_362 (.A(pwm_cnt[6]), .B(duty1[6]), 
         .Z(n38367)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i13_2_lut_rep_362.init = 16'h6666;
    FD1S3IX duty1_i11 (.D(duty1_14__N_458[11]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i11.GSR = "DISABLED";
    FD1S3IX duty1_i10 (.D(duty1_14__N_458[10]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i10.GSR = "DISABLED";
    LUT4 i31941_2_lut_3_lut_4_lut (.A(pwm_cnt[6]), .B(duty1[6]), .C(duty1[5]), 
         .D(pwm_cnt[5]), .Z(n36777)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i31941_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_13_i2276_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[6]), 
         .D(n3351_adj_1563), .Z(n13_adj_1564)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2276_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX duty1_i9 (.D(duty1_14__N_458[9]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i9.GSR = "DISABLED";
    LUT4 pwm_cnt_14__I_0_53_i10_3_lut_3_lut (.A(pwm_cnt[6]), .B(duty1[6]), 
         .C(duty1[5]), .Z(n10_adj_1565)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i10_3_lut_3_lut.init = 16'hd4d4;
    FD1S3JX duty1_i8 (.D(duty1_14__N_458[8]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i8.GSR = "DISABLED";
    FD1S3JX duty1_i7 (.D(duty1_14__N_458[7]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i7.GSR = "DISABLED";
    FD1S3IX duty1_i6 (.D(duty1_14__N_458[6]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i6.GSR = "DISABLED";
    FD1S3JX duty1_i5 (.D(duty1_14__N_458[5]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i5.GSR = "DISABLED";
    FD1S3IX duty1_i4 (.D(duty1_14__N_458[4]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i4.GSR = "DISABLED";
    FD1S3IX duty1_i3 (.D(duty1_14__N_458[3]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i3.GSR = "DISABLED";
    FD1S3JX duty1_i2 (.D(duty1_14__N_458[2]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i2.GSR = "DISABLED";
    FD1S3JX duty1_i1 (.D(duty1_14__N_458[1]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty1_i1.GSR = "DISABLED";
    FD1S3JX duty0_i14 (.D(duty0_14__N_410[14]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i14.GSR = "DISABLED";
    FD1S3JX duty0_i13 (.D(duty0_14__N_410[13]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i13.GSR = "DISABLED";
    FD1S3IX duty0_i12 (.D(duty0_14__N_410[12]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i12.GSR = "DISABLED";
    FD1S3IX duty0_i11 (.D(duty0_14__N_410[11]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i11.GSR = "DISABLED";
    FD1S3IX duty0_i10 (.D(duty0_14__N_410[10]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i10.GSR = "DISABLED";
    FD1S3IX duty0_i9 (.D(duty0_14__N_410[9]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i9.GSR = "DISABLED";
    FD1S3JX duty0_i8 (.D(duty0_14__N_410[8]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i8.GSR = "DISABLED";
    FD1S3JX duty0_i7 (.D(duty0_14__N_410[7]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i7.GSR = "DISABLED";
    FD1S3IX duty0_i6 (.D(duty0_14__N_410[6]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i6.GSR = "DISABLED";
    FD1S3JX duty0_i5 (.D(duty0_14__N_410[5]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i5.GSR = "DISABLED";
    FD1S3IX duty0_i4 (.D(duty0_14__N_410[4]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i4.GSR = "DISABLED";
    FD1S3IX duty0_i3 (.D(duty0_14__N_410[3]), .CK(fastclk_c), .CD(n12416), 
            .Q(duty0[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i3.GSR = "DISABLED";
    FD1S3JX duty0_i2 (.D(duty0_14__N_410[2]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i2.GSR = "DISABLED";
    FD1S3JX duty0_i1 (.D(duty0_14__N_410[1]), .CK(fastclk_c), .PD(n12416), 
            .Q(duty0[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(41[10] 89[6])
    defparam duty0_i1.GSR = "DISABLED";
    LUT4 div_13_i1919_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[28]), 
         .D(n2834_adj_640), .Z(n2933)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1919_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1043_7 (.A0(n1412[25]), .B0(n1511_adj_2191[25]), .C0(GND_net), 
          .D0(n38305), .A1(n38305), .B1(n1412[26]), .C1(n1511_adj_2191[26]), 
          .D1(GND_net), .CIN(n30620), .COUT(n30621), .S0(n1610_adj_2187[25]), 
          .S1(n1610_adj_2187[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_7.INIT0 = 16'h303f;
    defparam div_9_add_1043_7.INIT1 = 16'hf000;
    defparam div_9_add_1043_7.INJECT1_0 = "NO";
    defparam div_9_add_1043_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1043_5 (.A0(n38305), .B0(n1412[23]), .C0(n1511_adj_2191[23]), 
          .D0(GND_net), .A1(n38305), .B1(n1412[24]), .C1(n1511_adj_2191[24]), 
          .D1(GND_net), .CIN(n30619), .COUT(n30620), .S0(n1610_adj_2187[23]), 
          .S1(n1610_adj_2187[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_5.INIT0 = 16'hf000;
    defparam div_9_add_1043_5.INIT1 = 16'hf000;
    defparam div_9_add_1043_5.INJECT1_0 = "NO";
    defparam div_9_add_1043_5.INJECT1_1 = "NO";
    LUT4 div_13_i2258_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[24]), 
         .D(n3333_adj_1572), .Z(n49)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2258_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_842_Select_13_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[13]), 
         .D(n2983), .Z(duty0_14__N_410[13])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_13_i4_3_lut_4_lut.init = 16'hff10;
    LUT4 div_13_i2251_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3392_adj_2177[31]), 
         .D(n3326_adj_1574), .Z(n63_adj_1575)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2251_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1190_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[20]), 
         .D(n1753_adj_1268), .Z(n1852)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2412_3_lut_4_lut (.A(n28484), .B(n13621), .C(n3556), 
         .D(n4990[6]), .Z(n197[6])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2412_3_lut_4_lut.init = 16'hfe0e;
    LUT4 div_13_i2417_3_lut_4_lut (.A(n28267), .B(n13608), .C(n3556), 
         .D(n4990[1]), .Z(n197[1])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2417_3_lut_4_lut.init = 16'hfe0e;
    LUT4 div_13_i1922_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[25]), 
         .D(n2837), .Z(n2936_adj_1577)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1922_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1187_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[23]), 
         .D(n1750_adj_1073), .Z(n1849_adj_960)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1187_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1925_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[22]), 
         .D(n2840), .Z(n2939_adj_1579)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1925_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1192_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[18]), 
         .D(n333), .Z(n1854_adj_968)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_53_i15_2_lut_rep_363 (.A(pwm_cnt[7]), .B(duty1[7]), 
         .Z(n38368)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i15_2_lut_rep_363.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_53_i12_3_lut_3_lut (.A(pwm_cnt[7]), .B(duty1[7]), 
         .C(n10_adj_1565), .Z(n12_adj_1406)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i12_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_13_add_976_9 (.A0(n28420), .B0(n30262), .C0(n446), .D0(n1412_adj_2192[28]), 
          .A1(n28420), .B1(n30262), .C1(n446), .D1(n1412_adj_2192[29]), 
          .CIN(n30862), .COUT(n30863), .S0(n1511[28]), .S1(n1511[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_976_9.INIT0 = 16'hc0c0;
    defparam div_13_add_976_9.INIT1 = 16'h0000;
    defparam div_13_add_976_9.INJECT1_0 = "NO";
    defparam div_13_add_976_9.INJECT1_1 = "NO";
    LUT4 div_13_i1916_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[31]), 
         .D(n2831), .Z(n2930_adj_1583)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1916_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2253_3_lut_rep_164 (.A(n3328), .B(n3392_adj_2163[29]), 
         .C(n3359), .Z(n38169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2253_3_lut_rep_164.init = 16'hcaca;
    LUT4 div_13_i1939_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[8]), 
         .D(n2854_adj_601), .Z(n2953_adj_1586)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1939_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1191_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[19]), 
         .D(n1754_adj_1076), .Z(n1853_adj_967)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1188_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[22]), 
         .D(n1751_adj_1229), .Z(n1850_adj_964)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_157 (.A(n3328), .B(n3392_adj_2163[29]), .C(n3359), 
         .D(n38170), .Z(n34746)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_157.init = 16'hffca;
    LUT4 div_13_i1929_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[18]), 
         .D(n38227), .Z(n2943_adj_1588)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1929_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1931_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[16]), 
         .D(n2846_adj_615), .Z(n2945_adj_1590)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1931_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_then_3_lut (.A(n4540[23]), .B(n4540[3]), .C(n4540[5]), 
         .Z(n38417)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam i1_4_lut_then_3_lut.init = 16'hfefe;
    LUT4 div_13_i1928_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[19]), 
         .D(n2843_adj_637), .Z(n2942_adj_1592)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1928_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1713_17 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[25]), 
          .D0(n38266), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[26]), 
          .D1(n38265), .CIN(n30718), .COUT(n30719), .S0(n2600_adj_2186[25]), 
          .S1(n2600_adj_2186[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_17.INJECT1_0 = "NO";
    defparam div_9_add_1713_17.INJECT1_1 = "NO";
    CCU2C div_13_add_976_7 (.A0(n446), .B0(GND_net), .C0(n1412_adj_2192[26]), 
          .D0(n1351), .A1(n446), .B1(GND_net), .C1(n1412_adj_2192[27]), 
          .D1(n1350), .CIN(n30861), .COUT(n30862), .S0(n1511[26]), .S1(n1511[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_976_7.INIT0 = 16'h0c3f;
    defparam div_13_add_976_7.INIT1 = 16'hf3c0;
    defparam div_13_add_976_7.INJECT1_0 = "NO";
    defparam div_13_add_976_7.INJECT1_1 = "NO";
    CCU2C div_13_add_976_5 (.A0(n446), .B0(GND_net), .C0(n1412_adj_2192[24]), 
          .D0(n1353), .A1(n446), .B1(GND_net), .C1(n1412_adj_2192[25]), 
          .D1(n1352), .CIN(n30860), .COUT(n30861), .S0(n1511[24]), .S1(n1511[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_976_5.INIT0 = 16'hf3c0;
    defparam div_13_add_976_5.INIT1 = 16'hf3c0;
    defparam div_13_add_976_5.INJECT1_0 = "NO";
    defparam div_13_add_976_5.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i11_2_lut_rep_364 (.A(pwm_cnt[5]), .B(duty2[5]), 
         .Z(n38369)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i11_2_lut_rep_364.init = 16'h6666;
    LUT4 div_9_i1182_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[28]), 
         .D(n1745), .Z(n1844)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1182_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1713_15 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[23]), 
          .D0(n2443_adj_1319), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[24]), 
          .D1(n2442_adj_1601), .CIN(n30717), .COUT(n30718), .S0(n2600_adj_2186[23]), 
          .S1(n2600_adj_2186[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_15.INJECT1_0 = "NO";
    defparam div_9_add_1713_15.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i29_2_lut_rep_365 (.A(pwm_cnt[14]), .B(duty2[14]), 
         .Z(n38370)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i29_2_lut_rep_365.init = 16'h6666;
    CCU2C div_9_add_1713_13 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[21]), 
          .D0(n2445_adj_1311), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[22]), 
          .D1(n2444_adj_1604), .CIN(n30716), .COUT(n30717), .S0(n2600_adj_2186[21]), 
          .S1(n2600_adj_2186[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_13.INJECT1_0 = "NO";
    defparam div_9_add_1713_13.INJECT1_1 = "NO";
    LUT4 div_9_i1183_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[27]), 
         .D(n1746_adj_1208), .Z(n1845_adj_974)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1183_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1184_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[26]), 
         .D(n1747_adj_1206), .Z(n1846_adj_956)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_52_i14_3_lut_3_lut (.A(pwm_cnt[14]), .B(duty2[14]), 
         .C(duty2[13]), .Z(n14_adj_1341)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i14_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1713_11 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[19]), 
          .D0(n2447_adj_1320), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[20]), 
          .D1(n2446_adj_1313), .CIN(n30715), .COUT(n30716), .S0(n2600_adj_2186[19]), 
          .S1(n2600_adj_2186[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_11.INJECT1_0 = "NO";
    defparam div_9_add_1713_11.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i13_2_lut_rep_366 (.A(pwm_cnt[6]), .B(duty2[6]), 
         .Z(n38371)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i13_2_lut_rep_366.init = 16'h6666;
    LUT4 i31998_2_lut_3_lut_4_lut (.A(pwm_cnt[6]), .B(duty2[6]), .C(duty2[5]), 
         .D(pwm_cnt[5]), .Z(n36834)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i31998_2_lut_3_lut_4_lut.init = 16'h9009;
    CCU2C div_9_add_1713_9 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[17]), 
          .D0(n2449_adj_1322), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[18]), 
          .D1(n2448_adj_1321), .CIN(n30714), .COUT(n30715), .S0(n2600_adj_2186[17]), 
          .S1(n2600_adj_2186[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1713_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1713_9.INJECT1_0 = "NO";
    defparam div_9_add_1713_9.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i10_3_lut_3_lut (.A(pwm_cnt[6]), .B(duty2[6]), 
         .C(duty2[5]), .Z(n10_adj_1609)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i10_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_13_add_976_3 (.A0(n446), .B0(GND_net), .C0(n1412_adj_2192[22]), 
          .D0(n329), .A1(n446), .B1(GND_net), .C1(n1412_adj_2192[23]), 
          .D1(n1354), .CIN(n30859), .COUT(n30860), .S0(n1511[22]), .S1(n1511[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_976_3.INIT0 = 16'hf3c0;
    defparam div_13_add_976_3.INIT1 = 16'h0c3f;
    defparam div_13_add_976_3.INJECT1_0 = "NO";
    defparam div_13_add_976_3.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i15_2_lut_rep_367 (.A(pwm_cnt[7]), .B(duty2[7]), 
         .Z(n38372)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i15_2_lut_rep_367.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_52_i12_3_lut_3_lut (.A(pwm_cnt[7]), .B(duty2[7]), 
         .C(n10_adj_1609), .Z(n12_adj_1177)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i12_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1713_7 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[15]), 
          .D0(n2451_adj_1323), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[16]), 
          .D1(n2450_adj_1324), .CIN(n30713), .COUT(n30714), .S0(n2600_adj_2186[15]), 
          .S1(n2600_adj_2186[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1713_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1713_7.INJECT1_0 = "NO";
    defparam div_9_add_1713_7.INJECT1_1 = "NO";
    LUT4 rem_10_i2257_3_lut_rep_165 (.A(n3332), .B(n3392_adj_2163[25]), 
         .C(n3359), .Z(n38170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2257_3_lut_rep_165.init = 16'hcaca;
    LUT4 div_13_i1936_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[11]), 
         .D(n2851_adj_647), .Z(n2950_adj_1616)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1936_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_976_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n330), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30859), .S1(n1511[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_976_1.INIT0 = 16'h0000;
    defparam div_13_add_976_1.INIT1 = 16'h555a;
    defparam div_13_add_976_1.INJECT1_0 = "NO";
    defparam div_13_add_976_1.INJECT1_1 = "NO";
    LUT4 div_9_i1181_3_lut_4_lut (.A(n28287), .B(n13653), .C(n1808_adj_2179[29]), 
         .D(n1744_adj_520), .Z(n1843)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1181_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1924_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[23]), 
         .D(n2839_adj_643), .Z(n2938_adj_1618)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1924_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1933_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[14]), 
         .D(n2848_adj_646), .Z(n2947_adj_1620)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1933_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_158 (.A(n3332), .B(n3392_adj_2163[25]), .C(n3359), 
         .D(n3433), .Z(n35486)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_158.init = 16'hffca;
    LUT4 i1_4_lut_else_3_lut (.A(n13549), .B(n28574), .C(n13547), .D(n28588), 
         .Z(n38416)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam i1_4_lut_else_3_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_159 (.A(n2939), .B(n2996_adj_2193[22]), .C(n38217), 
         .D(n3044_adj_1296), .Z(n35142)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_159.init = 16'hffca;
    LUT4 rem_10_i2258_3_lut_rep_166 (.A(n3333), .B(n3392_adj_2163[24]), 
         .C(n3359), .Z(n38171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2258_3_lut_rep_166.init = 16'hcaca;
    LUT4 i28737_2_lut_rep_289 (.A(n1610[30]), .B(n28558), .Z(n38294)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i28737_2_lut_rep_289.init = 16'h8888;
    LUT4 select_842_Select_5_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[5]), 
         .D(n2983), .Z(duty0_14__N_410[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_5_i4_3_lut_4_lut.init = 16'hff10;
    LUT4 i1_2_lut_4_lut_adj_160 (.A(n3333), .B(n3392_adj_2163[24]), .C(n3359), 
         .D(n3433), .Z(n34740)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_160.init = 16'hffca;
    LUT4 i1_4_lut_4_lut (.A(n1610[30]), .B(n28558), .C(n33572), .D(n1646), 
         .Z(n13640)) /* synthesis lut_function=(A (B+(D))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_4_lut.init = 16'hffc8;
    LUT4 i24187_2_lut_rep_290 (.A(n28090), .B(n13631), .Z(n38295)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24187_2_lut_rep_290.init = 16'heeee;
    LUT4 rem_10_i1181_3_lut_rep_285_4_lut (.A(n28090), .B(n13631), .C(n1808[29]), 
         .D(n1744), .Z(n38290)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1181_3_lut_rep_285_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_161 (.A(n2953), .B(n2996_adj_2193[8]), .C(n38217), 
         .D(n3051_adj_1624), .Z(n34720)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_161.init = 16'hca00;
    LUT4 i24498_2_lut_rep_212 (.A(n28436), .B(n13592), .Z(n38217)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24498_2_lut_rep_212.init = 16'heeee;
    LUT4 rem_10_i1983_3_lut_rep_205_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[31]), 
         .D(n2930), .Z(n38210)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1983_3_lut_rep_205_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1992_3_lut_rep_210_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[22]), 
         .D(n2939), .Z(n38215)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1992_3_lut_rep_210_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_162 (.A(n3232_adj_766), .B(n3293_adj_2164[26]), 
         .C(n38176), .D(n3330_adj_613), .Z(n35302)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_162.init = 16'hffca;
    LUT4 rem_10_i2006_3_lut_rep_211_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[8]), 
         .D(n2953), .Z(n38216)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2006_3_lut_rep_211_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_163 (.A(n3238_adj_754), .B(n3293_adj_2164[20]), 
         .C(n38176), .D(n3341_adj_604), .Z(n35318)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_163.init = 16'hffca;
    LUT4 rem_10_i1985_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[29]), 
         .D(n2932), .Z(n3031_adj_1629)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1985_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_164 (.A(n3253_adj_657), .B(n3293_adj_2164[5]), 
         .C(n38176), .D(n3351_adj_1563), .Z(n34904)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_164.init = 16'hca00;
    LUT4 rem_10_i1998_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[16]), 
         .D(n2945), .Z(n3044_adj_1296)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1998_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1182_3_lut_rep_286_4_lut (.A(n28090), .B(n13631), .C(n1808[28]), 
         .D(n1745_adj_1502), .Z(n38291)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1182_3_lut_rep_286_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_909_11 (.A0(n38[28]), .B0(n3556), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n30858), 
          .S0(n1412_adj_2192[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_909_11.INIT0 = 16'hfff0;
    defparam div_13_add_909_11.INIT1 = 16'h0000;
    defparam div_13_add_909_11.INJECT1_0 = "NO";
    defparam div_13_add_909_11.INJECT1_1 = "NO";
    LUT4 rem_10_i1190_3_lut_rep_287_4_lut (.A(n28090), .B(n13631), .C(n1808[20]), 
         .D(n1753), .Z(n38292)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1190_3_lut_rep_287_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2342_3_lut_4_lut (.A(n3450), .B(n38178), .C(n3458), .D(n3449), 
         .Z(n3548)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2342_3_lut_4_lut.init = 16'h1fe0;
    LUT4 i24578_2_lut_rep_171 (.A(n28528), .B(n13610), .Z(n38176)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24578_2_lut_rep_171.init = 16'heeee;
    LUT4 pwm_cnt_14__I_0_51_i11_2_lut_rep_368 (.A(pwm_cnt[5]), .B(duty3[5]), 
         .Z(n38373)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i11_2_lut_rep_368.init = 16'h6666;
    LUT4 rem_10_i1999_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[15]), 
         .D(n2946), .Z(n3045_adj_1633)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1999_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1713_5 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[13]), 
          .D0(n2453_adj_1327), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[14]), 
          .D1(n2452_adj_1325), .CIN(n30712), .COUT(n30713), .S0(n2600_adj_2186[13]), 
          .S1(n2600_adj_2186[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1713_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1713_5.INJECT1_0 = "NO";
    defparam div_9_add_1713_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_175 (.A(n3352), .B(n3353_adj_1636), .C(n3354_adj_1637), 
         .Z(n38180)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_175.init = 16'h8080;
    LUT4 div_13_i1117_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[26]), 
         .D(n1351), .Z(n1747_adj_1430)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3397_bdd_4_lut_adj_165 (.A(n3327), .B(n3330), .C(n3340), .D(n3343), 
         .Z(n38058)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3397_bdd_4_lut_adj_165.init = 16'hfffe;
    LUT4 div_13_i2210_3_lut_rep_169_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[5]), 
         .D(n3253_adj_657), .Z(n38174)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2210_3_lut_rep_169_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1997_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[17]), 
         .D(n2944), .Z(n3043_adj_1639)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1997_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1179_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[31]), 
         .D(n1742_adj_1640), .Z(n1841)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1179_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1986_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[28]), 
         .D(n38220), .Z(n3032_adj_1642)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1986_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1180_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[30]), 
         .D(n1743_adj_1643), .Z(n1842)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2195_3_lut_rep_168_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[20]), 
         .D(n3238_adj_754), .Z(n38173)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2195_3_lut_rep_168_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1994_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[20]), 
         .D(n38225), .Z(n3040_adj_1645)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1994_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1192_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[18]), 
         .D(n582), .Z(n1854)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1186_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[24]), 
         .D(n1749), .Z(n1848)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1186_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1043_3 (.A0(n38307), .B0(n1511_adj_2191[21]), .C0(n35[19]), 
          .D0(GND_net), .A1(n1412[22]), .B1(n1511_adj_2191[22]), .C1(n38305), 
          .D1(GND_net), .CIN(n30618), .COUT(n30619), .S0(n1610_adj_2187[21]), 
          .S1(n1610_adj_2187[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_3.INIT0 = 16'hcca0;
    defparam div_9_add_1043_3.INIT1 = 16'h330f;
    defparam div_9_add_1043_3.INJECT1_0 = "NO";
    defparam div_9_add_1043_3.INJECT1_1 = "NO";
    LUT4 div_13_i2208_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[7]), 
         .D(n3251_adj_672), .Z(n3350_adj_1649)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2208_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2000_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[14]), 
         .D(n2947_adj_571), .Z(n3046_adj_1651)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2000_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1189_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[21]), 
         .D(n1752), .Z(n1851)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1189_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1996_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[18]), 
         .D(n2943), .Z(n3042_adj_1653)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1996_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2198_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[17]), 
         .D(n3241_adj_685), .Z(n3340_adj_1655)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2198_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1989_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[25]), 
         .D(n2936), .Z(n3035_adj_1657)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1989_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3397_bdd_4_lut_32455 (.A(n3392_adj_2163[27]), .B(n3392_adj_2163[30]), 
         .C(n3392_adj_2163[17]), .D(n3392_adj_2163[14]), .Z(n38057)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3397_bdd_4_lut_32455.init = 16'hfffe;
    LUT4 rem_10_i1187_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[23]), 
         .D(n1750), .Z(n1849)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1187_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1993_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[21]), 
         .D(n2940), .Z(n3039_adj_1663)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1993_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1984_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[30]), 
         .D(n2931_adj_535), .Z(n3030_adj_1665)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1984_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1188_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[22]), 
         .D(n1751), .Z(n1850)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1991_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[23]), 
         .D(n2938), .Z(n3037_adj_1667)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1991_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2196_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[19]), 
         .D(n3239_adj_773), .Z(n3338_adj_1307)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2196_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1987_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[27]), 
         .D(n2934), .Z(n3033_adj_1670)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1987_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2191_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[24]), 
         .D(n3234_adj_688), .Z(n3333_adj_1572)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3359_bdd_4_lut_32313 (.A(n3392[30]), .B(n3392[20]), .C(n3392[25]), 
         .D(n3392[14]), .Z(n37664)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3359_bdd_4_lut_32313.init = 16'hfffe;
    LUT4 rem_10_i1990_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[24]), 
         .D(n2937_adj_526), .Z(n3036_adj_1673)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1990_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1995_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[19]), 
         .D(n2942), .Z(n3041_adj_1675)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1995_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1184_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[26]), 
         .D(n1747), .Z(n1846)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2189_3_lut_rep_167_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[26]), 
         .D(n3232_adj_766), .Z(n38172)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2189_3_lut_rep_167_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_909_9 (.A0(n38[27]), .B0(n38298), .C0(n3556), .D0(n38[28]), 
          .A1(n38[28]), .B1(n3556), .C1(GND_net), .D1(VCC_net), .CIN(n30857), 
          .COUT(n30858), .S0(n1412_adj_2192[29]), .S1(n1412_adj_2192[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_909_9.INIT0 = 16'h0000;
    defparam div_13_add_909_9.INIT1 = 16'h0000;
    defparam div_13_add_909_9.INJECT1_0 = "NO";
    defparam div_13_add_909_9.INJECT1_1 = "NO";
    LUT4 div_9_i2128_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[20]), 
         .D(n3139), .Z(n3238)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2128_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1988_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[26]), 
         .D(n2935), .Z(n3034_adj_1677)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1988_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2007_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[7]), 
         .D(n2954), .Z(n3053_adj_1679)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2007_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_909_7 (.A0(n38298), .B0(n38[28]), .C0(n3556), .D0(n38[27]), 
          .A1(n38[27]), .B1(n38298), .C1(n3556), .D1(n38[28]), .CIN(n30856), 
          .COUT(n30857), .S0(n1412_adj_2192[27]), .S1(n1412_adj_2192[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_909_7.INIT0 = 16'h8f7f;
    defparam div_13_add_909_7.INIT1 = 16'h8000;
    defparam div_13_add_909_7.INJECT1_0 = "NO";
    defparam div_13_add_909_7.INJECT1_1 = "NO";
    CCU2C div_13_add_909_5 (.A0(n1352), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n1351), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30855), 
          .COUT(n30856), .S0(n1412_adj_2192[25]), .S1(n1412_adj_2192[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_909_5.INIT0 = 16'haaaa;
    defparam div_13_add_909_5.INIT1 = 16'haaaa;
    defparam div_13_add_909_5.INJECT1_0 = "NO";
    defparam div_13_add_909_5.INJECT1_1 = "NO";
    CCU2C div_13_add_909_3 (.A0(n38[28]), .B0(n38[23]), .C0(n3556), .D0(n72_adj_5), 
          .A1(n1353), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30854), 
          .COUT(n30855), .S0(n1412_adj_2192[23]), .S1(n1412_adj_2192[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_909_3.INIT0 = 16'h6f60;
    defparam div_13_add_909_3.INIT1 = 16'h555a;
    defparam div_13_add_909_3.INJECT1_0 = "NO";
    defparam div_13_add_909_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1191_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[19]), 
         .D(n1754), .Z(n1853)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1648_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[31]), 
         .D(n38254), .Z(n2534)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1648_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_909_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n329), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n30854), .S1(n1412_adj_2192[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_909_1.INIT0 = 16'h0000;
    defparam div_13_add_909_1.INIT1 = 16'h555a;
    defparam div_13_add_909_1.INJECT1_0 = "NO";
    defparam div_13_add_909_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_909_11 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), .CIN(n30852), 
          .S0(n1412_adj_2194[30]), .S1(n1412_adj_2194[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_909_11.INIT0 = 16'h0000;
    defparam rem_10_add_909_11.INIT1 = 16'hffff;
    defparam rem_10_add_909_11.INJECT1_0 = "NO";
    defparam rem_10_add_909_11.INJECT1_1 = "NO";
    LUT4 div_13_i2201_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[14]), 
         .D(n3244_adj_807), .Z(n3343_adj_1209)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2201_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_909_9 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), .CIN(n30851), 
          .COUT(n30852), .S0(n1412_adj_2194[28]), .S1(n1412_adj_2194[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_909_9.INIT0 = 16'h2000;
    defparam rem_10_add_909_9.INIT1 = 16'h0000;
    defparam rem_10_add_909_9.INJECT1_0 = "NO";
    defparam rem_10_add_909_9.INJECT1_1 = "NO";
    LUT4 rem_10_i1183_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[27]), 
         .D(n1746), .Z(n1845)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1183_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2008_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[6]), 
         .D(n594), .Z(n3054_adj_1686)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2008_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_909_7 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), .CIN(n30850), 
          .COUT(n30851), .S0(n1412_adj_2194[26]), .S1(n1412_adj_2194[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_909_7.INIT0 = 16'h0000;
    defparam rem_10_add_909_7.INIT1 = 16'hffff;
    defparam rem_10_add_909_7.INJECT1_0 = "NO";
    defparam rem_10_add_909_7.INJECT1_1 = "NO";
    LUT4 rem_10_i1185_3_lut_4_lut (.A(n28090), .B(n13631), .C(n1808[25]), 
         .D(n1748), .Z(n1847)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2001_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[13]), 
         .D(n2948), .Z(n3047_adj_1690)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2001_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1053_3_lut_rep_291 (.A(n1354), .B(n1610[23]), .C(n28558), 
         .Z(n38296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1053_3_lut_rep_291.init = 16'hcaca;
    LUT4 rem_10_i2002_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[12]), 
         .D(n2949), .Z(n3048_adj_1692)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2002_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_166 (.A(n1354), .B(n1610[23]), .C(n28558), 
         .D(n1652), .Z(n34782)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_166.init = 16'hca00;
    LUT4 rem_10_i2003_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[11]), 
         .D(n2950), .Z(n3049_adj_1694)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2003_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2185_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[30]), 
         .D(n3228_adj_682), .Z(n3327_adj_632)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2005_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[9]), 
         .D(n38224), .Z(n3051_adj_1624)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2005_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i848_3_lut_4_lut (.A(n38303), .B(n6_adj_1495), .C(n446), 
         .D(n38301), .Z(n1350)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i848_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_3_lut_4_lut (.A(n38301), .B(n38303), .C(n446), .D(n6_adj_1495), 
         .Z(n1448)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 div_13_i2192_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[23]), 
         .D(n3235_adj_792), .Z(n3334_adj_1561)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2187_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[28]), 
         .D(n38182), .Z(n3329)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2187_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2004_3_lut_4_lut (.A(n28436), .B(n13592), .C(n2996_adj_2193[10]), 
         .D(n2951), .Z(n3050_adj_1700)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2004_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4851_2_lut_rep_296 (.A(n38[27]), .B(n3556), .Z(n38301)) /* synthesis lut_function=(A (B)) */ ;
    defparam i4851_2_lut_rep_296.init = 16'h8888;
    LUT4 i24622_2_lut_rep_213 (.A(n28574), .B(n13549), .Z(n38218)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24622_2_lut_rep_213.init = 16'heeee;
    CCU2C div_9_add_1713_3 (.A0(n13554), .B0(n28319), .C0(n2501_adj_2190[11]), 
          .D0(n340_adj_1326), .A1(n13554), .B1(n28319), .C1(n2501_adj_2190[12]), 
          .D1(n2454_adj_1328), .CIN(n30711), .COUT(n30712), .S0(n2600_adj_2186[11]), 
          .S1(n2600_adj_2186[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1713_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1713_3.INJECT1_0 = "NO";
    defparam div_9_add_1713_3.INJECT1_1 = "NO";
    LUT4 div_9_i1984_3_lut_rep_207_4_lut (.A(n28574), .B(n13549), .C(n2996[30]), 
         .D(n2931), .Z(n38212)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1984_3_lut_rep_207_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_167 (.A(n38[27]), .B(n3556), .C(n6_adj_1495), 
         .D(n38303), .Z(n30262)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_167.init = 16'h8000;
    LUT4 div_9_i2005_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[9]), 
         .D(n2952), .Z(n3051)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2005_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1999_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[15]), 
         .D(n2946_adj_759), .Z(n3045)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1999_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i27_3_lut_rep_298 (.A(n63_adj_3), .B(n38[26]), .C(n3556), 
         .Z(n38303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i27_3_lut_rep_298.init = 16'hcaca;
    LUT4 i26256_2_lut_rep_293_4_lut (.A(n63_adj_3), .B(n38[26]), .C(n3556), 
         .D(n6_adj_1495), .Z(n38298)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i26256_2_lut_rep_293_4_lut.init = 16'hca00;
    LUT4 div_9_i2007_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[7]), 
         .D(n2954_adj_836), .Z(n3053)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2007_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2008_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[6]), 
         .D(n345), .Z(n3054)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2008_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2209_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[6]), 
         .D(n3252_adj_718), .Z(n3351_adj_1563)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2209_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1993_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[21]), 
         .D(n2940_adj_742), .Z(n3039)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1993_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_168 (.A(n3352), .B(n3353_adj_1636), .C(n3354_adj_1637), 
         .D(n3293[6]), .Z(n31_adj_1704)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_168.init = 16'hff80;
    LUT4 pwm_cnt_14__I_0_51_i29_2_lut_rep_369 (.A(pwm_cnt[14]), .B(duty3[14]), 
         .Z(n38374)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i29_2_lut_rep_369.init = 16'h6666;
    LUT4 div_9_i2003_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[11]), 
         .D(n2950_adj_820), .Z(n3049)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2003_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3409_bdd_4_lut_32319 (.A(n3392[15]), .B(n3392[22]), .C(n3392[23]), 
         .D(n3392[12]), .Z(n37670)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3409_bdd_4_lut_32319.init = 16'hfffe;
    LUT4 div_13_i1649_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[30]), 
         .D(n2436), .Z(n2535)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1649_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1659_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[20]), 
         .D(n2446), .Z(n2545)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1659_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1713_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[10]), .D1(duty0_14__N_426[8]), 
          .COUT(n30711), .S1(n2600_adj_2186[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1713_1.INIT0 = 16'h0000;
    defparam div_9_add_1713_1.INIT1 = 16'h04bf;
    defparam div_9_add_1713_1.INJECT1_0 = "NO";
    defparam div_9_add_1713_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1646_21 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[30]), 
          .D0(n2337_adj_1706), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[31]), 
          .D1(n2336_adj_1708), .CIN(n30709), .S0(n2501_adj_2190[30]), 
          .S1(n2501_adj_2190[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_21.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_21.INJECT1_0 = "NO";
    defparam div_9_add_1646_21.INJECT1_1 = "NO";
    LUT4 n3410_bdd_4_lut_32264 (.A(n3392_adj_2177[14]), .B(n3392_adj_2177[16]), 
         .C(n3392_adj_2177[18]), .D(n3392_adj_2177[10]), .Z(n37504)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3410_bdd_4_lut_32264.init = 16'hfffe;
    LUT4 n3409_bdd_4_lut (.A(n3342_adj_1713), .B(n3334_adj_1714), .C(n3345_adj_1715), 
         .D(n3335_adj_1716), .Z(n37671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3409_bdd_4_lut.init = 16'hfffe;
    LUT4 div_9_i2006_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[8]), 
         .D(n2953_adj_830), .Z(n3052)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2006_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1985_3_lut_rep_206_4_lut (.A(n28574), .B(n13549), .C(n2996[29]), 
         .D(n2932_adj_709), .Z(n38211)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1985_3_lut_rep_206_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1995_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[19]), 
         .D(n2942_adj_746), .Z(n3041)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1995_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1994_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[20]), 
         .D(n2941), .Z(n3040)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1994_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n3399_bdd_4_lut_32272 (.A(n3392_adj_2177[25]), .B(n3392_adj_2177[22]), 
         .C(n3392_adj_2177[30]), .D(n3392_adj_2177[12]), .Z(n37515)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3399_bdd_4_lut_32272.init = 16'hfffe;
    LUT4 div_13_i2200_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[15]), 
         .D(n3243_adj_692), .Z(n3342_adj_1516)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2200_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2212_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[3]), 
         .D(n348), .Z(n3354_adj_1637)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2212_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2004_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[10]), 
         .D(n2951_adj_819), .Z(n3050)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2004_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_169 (.A(n36078), .B(n36084), .C(n36074), .D(n36080), 
         .Z(n13547)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_169.init = 16'hfffe;
    LUT4 div_9_i2001_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[13]), 
         .D(n2948_adj_787), .Z(n3047)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2001_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2002_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[12]), 
         .D(n2949_adj_786), .Z(n3048)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2002_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2205_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[10]), 
         .D(n3248_adj_695), .Z(n3347_adj_1210)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2205_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1986_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[28]), 
         .D(n38221), .Z(n3032)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1986_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2207_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[8]), 
         .D(n3250_adj_704), .Z(n3349_adj_1724)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2207_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2204_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[11]), 
         .D(n3247_adj_811), .Z(n3346_adj_1509)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2204_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1996_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[18]), 
         .D(n2943_adj_745), .Z(n3042)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1996_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1988_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[26]), 
         .D(n2935_adj_710), .Z(n3034)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1988_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1987_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[27]), 
         .D(n2934_adj_711), .Z(n3033)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1987_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_170 (.A(n3144), .B(n3129), .C(n3137), .D(n3145), 
         .Z(n36078)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_170.init = 16'hfffe;
    LUT4 div_9_i2211_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[4]), 
         .D(n3254), .Z(n3353_adj_1636)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2211_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_171 (.A(n35[19]), .B(n38307), .C(n1709_adj_2160[24]), 
         .D(n1709_adj_2160[25]), .Z(n35834)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_171.init = 16'h8000;
    LUT4 div_13_i2194_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[21]), 
         .D(n3237_adj_662), .Z(n3336_adj_1521)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2194_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1991_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[23]), 
         .D(n2938_adj_741), .Z(n3037)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1991_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1666_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[13]), 
         .D(n2453), .Z(n2552)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1666_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1653_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[26]), 
         .D(n38255), .Z(n2539)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1653_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1997_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[17]), 
         .D(n2944_adj_748), .Z(n3043)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1997_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1998_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[16]), 
         .D(n2945_adj_747), .Z(n3044)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1998_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_172 (.A(n3131_adj_1727), .B(n36076), .C(n36056), 
         .D(n3146), .Z(n36084)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_172.init = 16'hfffe;
    LUT4 div_13_i1656_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[23]), 
         .D(n2443), .Z(n2542)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1656_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_173 (.A(n3136), .B(n3142), .C(n3132_adj_1728), .Z(n36074)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_3_lut_adj_173.init = 16'hfefe;
    LUT4 div_9_i1983_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[31]), 
         .D(n2930_adj_706), .Z(n3029)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1983_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_174 (.A(n3130), .B(n3141), .C(n3139), .D(n3140), 
         .Z(n36080)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_174.init = 16'hfffe;
    LUT4 div_13_i2186_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[29]), 
         .D(n3229_adj_723), .Z(n3328_adj_1306)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2186_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1043_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), 
          .COUT(n30618), .S1(n1610_adj_2187[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1043_1.INIT0 = 16'h0000;
    defparam div_9_add_1043_1.INIT1 = 16'hdfff;
    defparam div_9_add_1043_1.INJECT1_0 = "NO";
    defparam div_9_add_1043_1.INJECT1_1 = "NO";
    LUT4 div_9_i1992_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[22]), 
         .D(n2939_adj_740), .Z(n3038)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1992_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_175 (.A(n3138), .B(n3128_adj_1528), .C(n3134), .D(n3135), 
         .Z(n36076)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_175.init = 16'hfffe;
    CCU2C div_9_add_976_11 (.A0(n12154), .B0(n5), .C0(n35[19]), .D0(n1412[30]), 
          .A1(n12154), .B1(n5), .C1(n35[19]), .D1(n1412[31]), .CIN(n30616), 
          .S0(n1511_adj_2191[30]), .S1(n1511_adj_2191[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_976_11.INIT0 = 16'hffff;
    defparam div_9_add_976_11.INIT1 = 16'hffff;
    defparam div_9_add_976_11.INJECT1_0 = "NO";
    defparam div_9_add_976_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_176 (.A(n35780), .B(n28184), .C(n3150), .D(n38200), 
         .Z(n28588)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_176.init = 16'ha8a0;
    LUT4 div_9_i1989_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[25]), 
         .D(n2936_adj_737), .Z(n3035)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1989_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2188_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[27]), 
         .D(n3231), .Z(n3330_adj_812)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2193_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[22]), 
         .D(n3236_adj_675), .Z(n3335_adj_635)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2193_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2000_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[14]), 
         .D(n2947), .Z(n3046)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2000_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_177 (.A(n3147), .B(n3148), .C(n3149), .Z(n35780)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_177.init = 16'h8080;
    LUT4 div_9_i1990_3_lut_4_lut (.A(n28574), .B(n13549), .C(n2996[24]), 
         .D(n2937), .Z(n3036)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1990_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2211_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[4]), 
         .D(n3254_adj_668), .Z(n3353_adj_1558)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2211_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24232_3_lut (.A(n347), .B(n3153), .C(n3154), .Z(n28184)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24232_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_4_lut_adj_178 (.A(n2734), .B(n2798[29]), .C(n38228), 
         .D(n2839_adj_643), .Z(n35462)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_178.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_179 (.A(n2834), .B(n2897_adj_2162[28]), .C(n38226), 
         .D(n2937_adj_526), .Z(n35206)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_179.init = 16'hffca;
    LUT4 rem_10_i2363_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[10]), 
         .D(n3545), .Z(n36[10])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2363_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_180 (.A(n2834_adj_880), .B(n2897[28]), .C(n38223), 
         .D(n2942_adj_746), .Z(n36134)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_180.init = 16'hffca;
    LUT4 div_13_i2190_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[25]), 
         .D(n3233_adj_795), .Z(n3332_adj_633)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_181 (.A(n2739), .B(n2798[24]), .C(n38228), 
         .D(n2840), .Z(n35466)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_181.init = 16'hffca;
    LUT4 rem_10_mux_3_i8_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[7]), .D(duty0_14__N_426[5]), 
         .Z(n593)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1857_i13_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[14]), .D(duty0_14__N_426[12]), 
         .Z(n337)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1857_i15_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[16]), .D(duty0_14__N_426[14]), 
         .Z(n335)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 div_13_i2212_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[3]), 
         .D(n348_adj_1735), .Z(n3354_adj_1736)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2212_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2372_3_lut_4_lut (.A(n5), .B(n38331), .C(n3568[1]), .D(n3458), 
         .Z(n36[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_i2372_3_lut_4_lut.init = 16'hf780;
    LUT4 i24618_2_lut_rep_218 (.A(n28568), .B(n13550), .Z(n38223)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24618_2_lut_rep_218.init = 16'heeee;
    LUT4 i1_3_lut_adj_182 (.A(n3194[7]), .B(n3194[9]), .C(n3194[8]), .Z(n34474)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_182.init = 16'h8080;
    LUT4 div_9_i1927_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[20]), 
         .D(n2842_adj_764), .Z(n2941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1927_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2416_3_lut_4_lut (.A(n28492), .B(n13629), .C(n38307), 
         .D(n4540[2]), .Z(n89[2])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_9_i2416_3_lut_4_lut.init = 16'hfe0e;
    LUT4 div_13_i1660_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[19]), 
         .D(n2447), .Z(n2546)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1660_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1857_i4_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[5]), .D(duty0_14__N_426[3]), 
         .Z(n346)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i4_3_lut_4_lut.init = 16'hf780;
    CCU2C div_9_add_1646_19 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[28]), 
          .D0(n2339_adj_1739), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[29]), 
          .D1(n2338_adj_1741), .CIN(n30708), .COUT(n30709), .S0(n2501_adj_2190[28]), 
          .S1(n2501_adj_2190[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_19.INJECT1_0 = "NO";
    defparam div_9_add_1646_19.INJECT1_1 = "NO";
    LUT4 mux_1857_i1_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[2]), .D(duty0_14__N_426[0]), 
         .Z(n349_adj_1742)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_183 (.A(n3293[9]), .B(n31_adj_1704), .C(n3293[8]), 
         .D(n3293[7]), .Z(n34078)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_183.init = 16'h8000;
    CCU2C div_9_add_976_9 (.A0(n12154), .B0(n5), .C0(n35[19]), .D0(n1412[28]), 
          .A1(n12154), .B1(n5), .C1(n35[19]), .D1(n1412[29]), .CIN(n30615), 
          .COUT(n30616), .S0(n1511_adj_2191[28]), .S1(n1511_adj_2191[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_976_9.INIT0 = 16'h4040;
    defparam div_9_add_976_9.INIT1 = 16'h0000;
    defparam div_9_add_976_9.INJECT1_0 = "NO";
    defparam div_9_add_976_9.INJECT1_1 = "NO";
    CCU2C div_9_add_1646_17 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[26]), 
          .D0(n2341_adj_1744), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[27]), 
          .D1(n2340_adj_1746), .CIN(n30707), .COUT(n30708), .S0(n2501_adj_2190[26]), 
          .S1(n2501_adj_2190[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_17.INJECT1_0 = "NO";
    defparam div_9_add_1646_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_909_5 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), .CIN(n30849), 
          .COUT(n30850), .S0(n1412_adj_2194[24]), .S1(n1412_adj_2194[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_909_5.INIT0 = 16'hffff;
    defparam rem_10_add_909_5.INIT1 = 16'h2000;
    defparam rem_10_add_909_5.INJECT1_0 = "NO";
    defparam rem_10_add_909_5.INJECT1_1 = "NO";
    LUT4 div_9_i2198_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[17]), 
         .D(n3241_adj_532), .Z(n3340_adj_1749)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2198_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_184 (.A(n34), .B(n38180), .C(n3252), .Z(n37_adj_1750)) /* synthesis lut_function=(A (B+(C))) */ ;
    defparam i1_3_lut_adj_184.init = 16'ha8a8;
    LUT4 mux_1857_i11_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[12]), .D(duty0_14__N_426[10]), 
         .Z(n339_adj_1752)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_mux_3_i5_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[4]), .D(duty0_14__N_426[2]), 
         .Z(n596)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_adj_185 (.A(n3392_adj_2177[7]), .B(n3392_adj_2177[9]), 
         .C(n3392_adj_2177[8]), .Z(n34015)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_185.init = 16'h8080;
    LUT4 i1_3_lut_adj_186 (.A(n3350_adj_1649), .B(n3349_adj_1724), .C(n3348_adj_1757), 
         .Z(n34013)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_186.init = 16'h8080;
    LUT4 i1_4_lut_adj_187 (.A(n35976), .B(n38164), .C(n31386), .D(n36690), 
         .Z(n34594)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_187.init = 16'h0002;
    LUT4 rem_10_mux_3_i10_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[9]), 
         .D(duty0_14__N_426[7]), .Z(n591)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_mux_3_i13_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[12]), 
         .D(duty0_14__N_426[10]), .Z(n588)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_rep_159_4_lut (.A(n5), .B(n38331), .C(n38165), .D(n33490), 
         .Z(n38164)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i1_3_lut_rep_159_4_lut.init = 16'hff80;
    LUT4 rem_10_mux_3_i6_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[5]), .D(duty0_14__N_426[3]), 
         .Z(n595)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 div_9_i1936_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[11]), 
         .D(n2851_adj_951), .Z(n2950_adj_820)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1936_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1857_i10_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[11]), .D(duty0_14__N_426[9]), 
         .Z(n340_adj_1326)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 div_9_i1938_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[9]), 
         .D(n2853_adj_954), .Z(n2952)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1938_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1932_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[15]), 
         .D(n2847_adj_934), .Z(n2946_adj_759)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1932_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1857_i2_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[3]), .D(duty0_14__N_426[1]), 
         .Z(n348)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i2_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_mux_3_i18_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[17]), 
         .D(duty0_14__N_426[15]), .Z(n583)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_1857_i3_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[4]), .D(duty0_14__N_426[2]), 
         .Z(n347)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_mux_3_i4_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[3]), .D(duty0_14__N_426[1]), 
         .Z(n597)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 rem_10_mux_3_i11_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[10]), 
         .D(duty0_14__N_426[8]), .Z(n590)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 div_9_i1939_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[8]), 
         .D(n2854_adj_955), .Z(n2953_adj_830)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1939_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_mux_3_i12_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[11]), 
         .D(duty0_14__N_426[9]), .Z(n589)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 div_13_i2206_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[9]), 
         .D(n3249_adj_698), .Z(n3348_adj_1757)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2206_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_mux_3_i17_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[16]), 
         .D(duty0_14__N_426[14]), .Z(n584)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 pwm_cnt_14__I_0_51_i14_3_lut_3_lut (.A(pwm_cnt[14]), .B(duty3[14]), 
         .C(duty3[13]), .Z(n14_adj_1343)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i14_3_lut_3_lut.init = 16'hd4d4;
    LUT4 rem_10_mux_3_i3_3_lut_4_lut (.A(n5), .B(n38331), .C(n2[2]), .D(duty0_14__N_426[0]), 
         .Z(n598)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam rem_10_mux_3_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_4_lut_adj_188 (.A(n3232_adj_1767), .B(n3293_adj_2161[26]), 
         .C(n38188), .D(n3335), .Z(n34818)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_188.init = 16'hffca;
    LUT4 pwm_cnt_14__I_0_51_i13_2_lut_rep_370 (.A(pwm_cnt[6]), .B(duty3[6]), 
         .Z(n38375)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i13_2_lut_rep_370.init = 16'h6666;
    LUT4 i32055_2_lut_3_lut_4_lut (.A(pwm_cnt[6]), .B(duty3[6]), .C(duty3[5]), 
         .D(pwm_cnt[5]), .Z(n36891)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32055_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 div_9_i1940_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[7]), 
         .D(n344), .Z(n2954_adj_836)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1940_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1646_15 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[24]), 
          .D0(n2343), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[25]), 
          .D1(n2342_adj_1771), .CIN(n30706), .COUT(n30707), .S0(n2501_adj_2190[24]), 
          .S1(n2501_adj_2190[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_15.INJECT1_0 = "NO";
    defparam div_9_add_1646_15.INJECT1_1 = "NO";
    LUT4 mux_1857_i8_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[9]), .D(duty0_14__N_426[7]), 
         .Z(n342_adj_1184)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 pwm_cnt_14__I_0_51_i10_3_lut_3_lut (.A(pwm_cnt[6]), .B(duty3[6]), 
         .C(duty3[5]), .Z(n10_adj_1772)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i10_3_lut_3_lut.init = 16'hd4d4;
    CCU2C rem_10_add_909_3 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), .CIN(n30848), 
          .COUT(n30849), .S0(n1412_adj_2194[22]), .S1(n1412_adj_2194[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_909_3.INIT0 = 16'h2000;
    defparam rem_10_add_909_3.INIT1 = 16'h0000;
    defparam rem_10_add_909_3.INJECT1_0 = "NO";
    defparam rem_10_add_909_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_909_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), 
          .COUT(n30848));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_909_1.INIT0 = 16'h000F;
    defparam rem_10_add_909_1.INIT1 = 16'hdfff;
    defparam rem_10_add_909_1.INJECT1_0 = "NO";
    defparam rem_10_add_909_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_976_13 (.A0(n12154), .B0(n5), .C0(n2[19]), .D0(n1412_adj_2194[31]), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n30847), 
          .S0(n1511_adj_2196[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_13.INIT0 = 16'hffff;
    defparam rem_10_add_976_13.INIT1 = 16'h0000;
    defparam rem_10_add_976_13.INJECT1_0 = "NO";
    defparam rem_10_add_976_13.INJECT1_1 = "NO";
    LUT4 div_13_i1665_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[14]), 
         .D(n2452), .Z(n2551)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1665_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1928_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[19]), 
         .D(n2843_adj_903), .Z(n2942_adj_746)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1928_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1251_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[26]), 
         .D(n1846_adj_1384), .Z(n1945_adj_1119)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1251_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_51_i15_2_lut_rep_371 (.A(pwm_cnt[7]), .B(duty3[7]), 
         .Z(n38376)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i15_2_lut_rep_371.init = 16'h6666;
    LUT4 div_9_i1937_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[10]), 
         .D(n2852_adj_953), .Z(n2951_adj_819)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1937_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i26533_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[26]), 
         .D(n35[19]), .Z(n1747_adj_1206)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26533_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1919_3_lut_rep_216_4_lut (.A(n28568), .B(n13550), .C(n2897[28]), 
         .D(n2834_adj_880), .Z(n38221)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1919_3_lut_rep_216_4_lut.init = 16'hf1e0;
    LUT4 i26530_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[30]), 
         .D(n35[19]), .Z(n1743)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26530_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26549_2_lut_rep_292_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[25]), 
         .D(n35[19]), .Z(n38297)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26549_2_lut_rep_292_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_189 (.A(n3253_adj_1776), .B(n3293_adj_2161[5]), 
         .C(n38188), .D(n3351), .Z(n34872)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_189.init = 16'hca00;
    LUT4 i26529_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[31]), 
         .D(n35[19]), .Z(n1742)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26529_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26532_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[27]), 
         .D(n35[19]), .Z(n1746_adj_1208)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26532_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26550_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[22]), 
         .D(n35[19]), .Z(n1751_adj_1229)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26550_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26535_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[23]), 
         .D(n35[19]), .Z(n1750_adj_1073)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26535_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26552_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[20]), 
         .D(n35[19]), .Z(n1753_adj_1268)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26552_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i24546_2_lut_rep_183 (.A(n28434), .B(n13620), .Z(n38188)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24546_2_lut_rep_183.init = 16'heeee;
    LUT4 i26548_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[28]), 
         .D(n35[19]), .Z(n1745)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26548_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 rem_10_i2187_3_lut_rep_179_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[28]), 
         .D(n3230_adj_1779), .Z(n38184)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2187_3_lut_rep_179_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1926_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[21]), 
         .D(n38236), .Z(n2940_adj_742)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1926_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1918_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[29]), 
         .D(n38230), .Z(n2932_adj_709)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1918_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_976_11 (.A0(n12154), .B0(n5), .C0(n2[19]), .D0(n1412_adj_2194[29]), 
          .A1(n12154), .B1(n5), .C1(n2[19]), .D1(n1412_adj_2194[30]), 
          .CIN(n30846), .COUT(n30847), .S0(n1511_adj_2196[29]), .S1(n1511_adj_2196[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_11.INIT0 = 16'h0000;
    defparam rem_10_add_976_11.INIT1 = 16'hffff;
    defparam rem_10_add_976_11.INJECT1_0 = "NO";
    defparam rem_10_add_976_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_976_9 (.A0(n12154), .B0(n5), .C0(n2[19]), .D0(n1412_adj_2194[27]), 
          .A1(n12154), .B1(n5), .C1(n2[19]), .D1(n1412_adj_2194[28]), 
          .CIN(n30845), .COUT(n30846), .S0(n1511_adj_2196[27]), .S1(n1511_adj_2196[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_9.INIT0 = 16'h0000;
    defparam rem_10_add_976_9.INIT1 = 16'h4040;
    defparam rem_10_add_976_9.INJECT1_0 = "NO";
    defparam rem_10_add_976_9.INJECT1_1 = "NO";
    LUT4 div_9_i1929_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[18]), 
         .D(n2844_adj_919), .Z(n2943_adj_745)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1929_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2184_3_lut_4_lut (.A(n28528), .B(n13610), .C(n3293_adj_2164[31]), 
         .D(n3227_adj_726), .Z(n3326_adj_1574)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2184_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1512_19 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[30]), 
          .D0(n2139_adj_1785), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[31]), 
          .D1(n2138_adj_1786), .CIN(n31270), .S0(n2303_adj_2197[30]), 
          .S1(n2303_adj_2197[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1512_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1512_19.INJECT1_0 = "NO";
    defparam rem_10_add_1512_19.INJECT1_1 = "NO";
    CCU2C rem_10_add_1512_17 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[28]), 
          .D0(n2141_adj_1789), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[29]), 
          .D1(n2140_adj_1790), .CIN(n31269), .COUT(n31270), .S0(n2303_adj_2197[28]), 
          .S1(n2303_adj_2197[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1512_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1512_17.INJECT1_0 = "NO";
    defparam rem_10_add_1512_17.INJECT1_1 = "NO";
    LUT4 i26534_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[24]), 
         .D(n35[19]), .Z(n1749_adj_1212)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26534_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26553_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[19]), 
         .D(n35[19]), .Z(n1754_adj_1076)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26553_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26551_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709_adj_2160[21]), 
         .D(n35[19]), .Z(n1752_adj_1270)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26551_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1935_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[12]), 
         .D(n2850_adj_952), .Z(n2949_adj_786)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1935_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1916_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[31]), 
         .D(n2831_adj_857), .Z(n2930_adj_706)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1916_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_976_7 (.A0(n12154), .B0(n5), .C0(n35[19]), .D0(n1412[26]), 
          .A1(n12154), .B1(n5), .C1(n35[19]), .D1(n1412[27]), .CIN(n30614), 
          .COUT(n30615), .S0(n1511_adj_2191[26]), .S1(n1511_adj_2191[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_976_7.INIT0 = 16'hffff;
    defparam div_9_add_976_7.INIT1 = 16'h0000;
    defparam div_9_add_976_7.INJECT1_0 = "NO";
    defparam div_9_add_976_7.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_51_i12_3_lut_3_lut (.A(pwm_cnt[7]), .B(duty3[7]), 
         .C(n10_adj_1772), .Z(n12_adj_841)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i12_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_9_i2118_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[30]), 
         .D(n3129), .Z(n3228)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2138_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[10]), 
         .D(n3149), .Z(n3248)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2138_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1921_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[26]), 
         .D(n2836_adj_888), .Z(n2935_adj_710)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1921_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1512_15 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[26]), 
          .D0(n2143_adj_1793), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[27]), 
          .D1(n2142_adj_1794), .CIN(n31268), .COUT(n31269), .S0(n2303_adj_2197[26]), 
          .S1(n2303_adj_2197[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1512_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1512_15.INJECT1_0 = "NO";
    defparam rem_10_add_1512_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_1512_13 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[24]), 
          .D0(n2145_adj_1797), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[25]), 
          .D1(n2144_adj_1798), .CIN(n31267), .COUT(n31268), .S0(n2303_adj_2197[24]), 
          .S1(n2303_adj_2197[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1512_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1512_13.INJECT1_0 = "NO";
    defparam rem_10_add_1512_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_976_7 (.A0(n12154), .B0(n5), .C0(n2[19]), .D0(n1412_adj_2194[25]), 
          .A1(n12154), .B1(n5), .C1(n2[19]), .D1(n1412_adj_2194[26]), 
          .CIN(n30844), .COUT(n30845), .S0(n1511_adj_2196[25]), .S1(n1511_adj_2196[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_7.INIT0 = 16'h4040;
    defparam rem_10_add_976_7.INIT1 = 16'hffff;
    defparam rem_10_add_976_7.INJECT1_0 = "NO";
    defparam rem_10_add_976_7.INJECT1_1 = "NO";
    CCU2C rem_10_add_1512_11 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[22]), 
          .D0(n2147_adj_1803), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[23]), 
          .D1(n2146_adj_1804), .CIN(n31266), .COUT(n31267), .S0(n2303_adj_2197[22]), 
          .S1(n2303_adj_2197[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1512_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1512_11.INJECT1_0 = "NO";
    defparam rem_10_add_1512_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1512_9 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[20]), 
          .D0(n2149_adj_1807), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[21]), 
          .D1(n2148_adj_1808), .CIN(n31265), .COUT(n31266), .S0(n2303_adj_2197[20]), 
          .S1(n2303_adj_2197[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1512_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1512_9.INJECT1_0 = "NO";
    defparam rem_10_add_1512_9.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i9_2_lut_rep_372 (.A(pwm_cnt[4]), .B(duty0[4]), 
         .Z(n38377)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i9_2_lut_rep_372.init = 16'h6666;
    LUT4 div_9_i1930_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[17]), 
         .D(n2845_adj_917), .Z(n2944_adj_748)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1930_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1646_13 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[22]), 
          .D0(n2345_adj_1812), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[23]), 
          .D1(n2344_adj_1814), .CIN(n30705), .COUT(n30706), .S0(n2501_adj_2190[22]), 
          .S1(n2501_adj_2190[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_13.INJECT1_0 = "NO";
    defparam div_9_add_1646_13.INJECT1_1 = "NO";
    LUT4 i26571_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[31]), 
         .D(n2[19]), .Z(n1742_adj_1640)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26571_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2C rem_10_add_1512_7 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[18]), 
          .D0(n2151_adj_1815), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[19]), 
          .D1(n2150_adj_1816), .CIN(n31264), .COUT(n31265), .S0(n2303_adj_2197[18]), 
          .S1(n2303_adj_2197[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1512_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1512_7.INJECT1_0 = "NO";
    defparam rem_10_add_1512_7.INJECT1_1 = "NO";
    CCU2C rem_10_add_1512_5 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[16]), 
          .D0(n2153_adj_1819), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[17]), 
          .D1(n2152_adj_1820), .CIN(n31263), .COUT(n31264), .S0(n2303_adj_2197[16]), 
          .S1(n2303_adj_2197[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1512_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1512_5.INJECT1_0 = "NO";
    defparam rem_10_add_1512_5.INJECT1_1 = "NO";
    LUT4 rem_10_i2189_3_lut_rep_181_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[26]), 
         .D(n3232_adj_1767), .Z(n38186)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2189_3_lut_rep_181_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1920_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[27]), 
         .D(n38231), .Z(n2934_adj_711)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1920_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32168_4_lut (.A(n36698), .B(n36660), .C(n36628), .D(n36630), 
         .Z(n14116)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam i32168_4_lut.init = 16'h0008;
    LUT4 i26537_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[23]), 
         .D(n2[19]), .Z(n1750)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26537_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1924_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[23]), 
         .D(n2839_adj_665), .Z(n2938_adj_741)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1924_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1934_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[13]), 
         .D(n2849_adj_939), .Z(n2948_adj_787)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1934_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i31862_4_lut (.A(pwm_cnt[5]), .B(n36656), .C(n36658), .D(pwm_cnt[14]), 
         .Z(n36698)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i31862_4_lut.init = 16'h8000;
    LUT4 i26558_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[20]), 
         .D(n2[19]), .Z(n1753)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26558_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1931_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[16]), 
         .D(n2846_adj_936), .Z(n2945_adj_747)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1931_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2412_3_lut_4_lut (.A(n28568), .B(n13550), .C(n38307), 
         .D(n4540[6]), .Z(n89[6])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_9_i2412_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i26564_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[25]), 
         .D(n2[19]), .Z(n1748)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26564_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2C rem_10_add_1512_3 (.A0(n13597), .B0(n28387), .C0(n2204_adj_2172[14]), 
          .D0(n586), .A1(n13597), .B1(n28387), .C1(n2204_adj_2172[15]), 
          .D1(n2154_adj_1823), .CIN(n31262), .COUT(n31263), .S0(n2303_adj_2197[14]), 
          .S1(n2303_adj_2197[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1512_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1512_3.INJECT1_0 = "NO";
    defparam rem_10_add_1512_3.INJECT1_1 = "NO";
    LUT4 i31827_2_lut (.A(pwm_cnt[13]), .B(pwm_cnt[1]), .Z(n36660)) /* synthesis lut_function=(A (B)) */ ;
    defparam i31827_2_lut.init = 16'h8888;
    LUT4 i26560_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[21]), 
         .D(n2[19]), .Z(n1752)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26560_2_lut_3_lut_4_lut.init = 16'h8000;
    CCU2C rem_10_add_1512_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n51), .D1(n2[13]), 
          .COUT(n31262), .S1(n2303_adj_2197[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1512_1.INIT0 = 16'h0000;
    defparam rem_10_add_1512_1.INIT1 = 16'habef;
    defparam rem_10_add_1512_1.INJECT1_0 = "NO";
    defparam rem_10_add_1512_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1579_21 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[31]), 
          .D0(n2237_adj_1827), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31261), .S0(n2402_adj_2198[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_21.INIT1 = 16'h0000;
    defparam rem_10_add_1579_21.INJECT1_0 = "NO";
    defparam rem_10_add_1579_21.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_190 (.A(pwm_cnt[6]), .B(pwm_cnt[10]), .C(pwm_cnt[12]), 
         .Z(n36628)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_190.init = 16'hfefe;
    CCU2C div_9_add_1646_11 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[20]), 
          .D0(n2347_adj_1830), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[21]), 
          .D1(n38270), .CIN(n30704), .COUT(n30705), .S0(n2501_adj_2190[20]), 
          .S1(n2501_adj_2190[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_11.INJECT1_0 = "NO";
    defparam div_9_add_1646_11.INJECT1_1 = "NO";
    LUT4 i26562_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[22]), 
         .D(n2[19]), .Z(n1751)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26562_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26556_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[19]), 
         .D(n2[19]), .Z(n1754)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26556_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26538_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[24]), 
         .D(n2[19]), .Z(n1749)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26538_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 div_9_i1925_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[22]), 
         .D(n2840_adj_899), .Z(n2939_adj_740)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1925_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i26565_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[26]), 
         .D(n2[19]), .Z(n1747)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26565_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26570_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[30]), 
         .D(n2[19]), .Z(n1743_adj_1643)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26570_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_191 (.A(pwm_cnt[9]), .B(pwm_cnt[4]), .C(pwm_cnt[11]), 
         .D(pwm_cnt[3]), .Z(n36630)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_191.init = 16'hfffe;
    LUT4 i31823_2_lut (.A(pwm_cnt[0]), .B(pwm_cnt[7]), .Z(n36656)) /* synthesis lut_function=(A (B)) */ ;
    defparam i31823_2_lut.init = 16'h8888;
    LUT4 i31825_2_lut (.A(pwm_cnt[8]), .B(pwm_cnt[2]), .Z(n36658)) /* synthesis lut_function=(A (B)) */ ;
    defparam i31825_2_lut.init = 16'h8888;
    LUT4 div_9_i1922_3_lut_4_lut (.A(n28568), .B(n13550), .C(n2897[25]), 
         .D(n2837_adj_886), .Z(n2936_adj_737)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1922_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1654_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[25]), 
         .D(n2441), .Z(n2540)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1654_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1579_19 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[29]), 
          .D0(n2239_adj_1832), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[30]), 
          .D1(n2238_adj_1833), .CIN(n31260), .COUT(n31261), .S0(n2402_adj_2198[29]), 
          .S1(n2402_adj_2198[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1579_19.INJECT1_0 = "NO";
    defparam rem_10_add_1579_19.INJECT1_1 = "NO";
    LUT4 div_9_i2142_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[6]), 
         .D(n3153), .Z(n3252)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2142_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1579_17 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[27]), 
          .D0(n2241_adj_1836), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[28]), 
          .D1(n2240_adj_1837), .CIN(n31259), .COUT(n31260), .S0(n2402_adj_2198[27]), 
          .S1(n2402_adj_2198[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1579_17.INJECT1_0 = "NO";
    defparam rem_10_add_1579_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_1579_15 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[25]), 
          .D0(n2243_adj_1840), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[26]), 
          .D1(n2242_adj_1841), .CIN(n31258), .COUT(n31259), .S0(n2402_adj_2198[25]), 
          .S1(n2402_adj_2198[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1579_15.INJECT1_0 = "NO";
    defparam rem_10_add_1579_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_1579_13 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[23]), 
          .D0(n2245_adj_1844), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[24]), 
          .D1(n2244_adj_1845), .CIN(n31257), .COUT(n31258), .S0(n2402_adj_2198[23]), 
          .S1(n2402_adj_2198[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1579_13.INJECT1_0 = "NO";
    defparam rem_10_add_1579_13.INJECT1_1 = "NO";
    LUT4 div_13_i1651_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[28]), 
         .D(n2438), .Z(n2537)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1651_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1579_11 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[21]), 
          .D0(n2247_adj_1848), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[22]), 
          .D1(n2246_adj_1849), .CIN(n31256), .COUT(n31257), .S0(n2402_adj_2198[21]), 
          .S1(n2402_adj_2198[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1579_11.INJECT1_0 = "NO";
    defparam rem_10_add_1579_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1579_9 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[19]), 
          .D0(n2249_adj_1852), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[20]), 
          .D1(n2248_adj_1853), .CIN(n31255), .COUT(n31256), .S0(n2402_adj_2198[19]), 
          .S1(n2402_adj_2198[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1579_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1579_9.INJECT1_0 = "NO";
    defparam rem_10_add_1579_9.INJECT1_1 = "NO";
    LUT4 div_13_i1668_3_lut_4_lut (.A(n28446), .B(n13627), .C(n2501[11]), 
         .D(n340), .Z(n2554)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1668_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1579_7 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[17]), 
          .D0(n2251_adj_1856), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[18]), 
          .D1(n2250_adj_1857), .CIN(n31254), .COUT(n31255), .S0(n2402_adj_2198[17]), 
          .S1(n2402_adj_2198[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1579_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1579_7.INJECT1_0 = "NO";
    defparam rem_10_add_1579_7.INJECT1_1 = "NO";
    CCU2C div_9_add_1646_9 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[18]), 
          .D0(n2349_adj_1861), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[19]), 
          .D1(n2348_adj_1863), .CIN(n30703), .COUT(n30704), .S0(n2501_adj_2190[18]), 
          .S1(n2501_adj_2190[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1646_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1646_9.INJECT1_0 = "NO";
    defparam div_9_add_1646_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_976_5 (.A0(n12154), .B0(n5), .C0(n2[19]), .D0(n1412_adj_2194[23]), 
          .A1(n12154), .B1(n5), .C1(n2[19]), .D1(n1412_adj_2194[24]), 
          .CIN(n30843), .COUT(n30844), .S0(n1511_adj_2196[23]), .S1(n1511_adj_2196[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_5.INIT0 = 16'hffff;
    defparam rem_10_add_976_5.INIT1 = 16'h0000;
    defparam rem_10_add_976_5.INJECT1_0 = "NO";
    defparam rem_10_add_976_5.INJECT1_1 = "NO";
    LUT4 rem_10_i2210_3_lut_rep_182_4_lut (.A(n28434), .B(n13620), .C(n3293_adj_2161[5]), 
         .D(n3253_adj_1776), .Z(n38187)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2210_3_lut_rep_182_4_lut.init = 16'hf1e0;
    LUT4 i26568_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[28]), 
         .D(n2[19]), .Z(n1745_adj_1502)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26568_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i26569_2_lut_3_lut_4_lut (.A(n5), .B(n38331), .C(n1709[29]), 
         .D(n2[19]), .Z(n1744)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam i26569_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_1857_i14_3_lut_4_lut (.A(n5), .B(n38331), .C(n35[15]), .D(duty0_14__N_426[13]), 
         .Z(n336)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(52[16] 56[10])
    defparam mux_1857_i14_3_lut_4_lut.init = 16'hf780;
    CCU2C div_9_add_976_5 (.A0(n12154), .B0(n5), .C0(n35[19]), .D0(n1412[24]), 
          .A1(n12154), .B1(n5), .C1(n35[19]), .D1(n1412[25]), .CIN(n30613), 
          .COUT(n30614), .S0(n1511_adj_2191[24]), .S1(n1511_adj_2191[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_976_5.INIT0 = 16'h0000;
    defparam div_9_add_976_5.INIT1 = 16'h4040;
    defparam div_9_add_976_5.INJECT1_0 = "NO";
    defparam div_9_add_976_5.INJECT1_1 = "NO";
    LUT4 i31902_3_lut_4_lut (.A(pwm_cnt[4]), .B(duty0[4]), .C(n38381), 
         .D(n38382), .Z(n36738)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i31902_3_lut_4_lut.init = 16'h0009;
    LUT4 div_13_i2408_3_lut_4_lut (.A(n28446), .B(n13627), .C(n3556), 
         .D(n4990[10]), .Z(n197[10])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2408_3_lut_4_lut.init = 16'hfe0e;
    CCU2C div_9_add_1646_7 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[16]), 
          .D0(n2351_adj_1867), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[17]), 
          .D1(n2350_adj_1869), .CIN(n30702), .COUT(n30703), .S0(n2501_adj_2190[16]), 
          .S1(n2501_adj_2190[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1646_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1646_7.INJECT1_0 = "NO";
    defparam div_9_add_1646_7.INJECT1_1 = "NO";
    LUT4 i24141_2_lut_rep_246 (.A(n28082), .B(n13601), .Z(n38251)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24141_2_lut_rep_246.init = 16'heeee;
    CCU2C rem_10_add_976_3 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n12154), .B1(n5), .C1(n2[19]), .D1(n1412_adj_2194[22]), 
          .CIN(n30842), .COUT(n30843), .S0(n1511_adj_2196[21]), .S1(n1511_adj_2196[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_3.INIT0 = 16'h2000;
    defparam rem_10_add_976_3.INIT1 = 16'h4040;
    defparam rem_10_add_976_3.INJECT1_0 = "NO";
    defparam rem_10_add_976_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1718_3_lut_rep_245_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[28]), 
         .D(n2537_adj_1498), .Z(n38250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1718_3_lut_rep_245_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_54_i21_2_lut_rep_373 (.A(pwm_cnt[10]), .B(duty0[10]), 
         .Z(n38378)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i21_2_lut_rep_373.init = 16'h6666;
    LUT4 div_9_i2129_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[19]), 
         .D(n3140), .Z(n3239)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2129_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_54_i23_2_lut_rep_374 (.A(pwm_cnt[11]), .B(duty0[11]), 
         .Z(n38379)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i23_2_lut_rep_374.init = 16'h6666;
    CCU2C rem_10_add_1579_5 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[15]), 
          .D0(n2253_adj_1872), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[16]), 
          .D1(n2252_adj_1873), .CIN(n31253), .COUT(n31254), .S0(n2402_adj_2198[15]), 
          .S1(n2402_adj_2198[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1579_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1579_5.INJECT1_0 = "NO";
    defparam rem_10_add_1579_5.INJECT1_1 = "NO";
    LUT4 i31911_2_lut_3_lut_4_lut (.A(pwm_cnt[11]), .B(duty0[11]), .C(duty0[10]), 
         .D(pwm_cnt[10]), .Z(n36747)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i31911_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 pwm_cnt_14__I_0_54_i18_3_lut_3_lut (.A(pwm_cnt[11]), .B(duty0[11]), 
         .C(duty0[10]), .Z(n18_adj_1876)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i18_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1646_5 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[14]), 
          .D0(n2353_adj_1878), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[15]), 
          .D1(n2352_adj_1880), .CIN(n30701), .COUT(n30702), .S0(n2501_adj_2190[14]), 
          .S1(n2501_adj_2190[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1646_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1646_5.INJECT1_0 = "NO";
    defparam div_9_add_1646_5.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i25_2_lut_rep_375 (.A(pwm_cnt[12]), .B(duty0[12]), 
         .Z(n38380)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i25_2_lut_rep_375.init = 16'h6666;
    CCU2C rem_10_add_976_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), 
          .COUT(n30842));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_976_1.INIT0 = 16'h000F;
    defparam rem_10_add_976_1.INIT1 = 16'hdfff;
    defparam rem_10_add_976_1.INJECT1_0 = "NO";
    defparam rem_10_add_976_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1043_13 (.A0(n38306), .B0(n1412_adj_2194[30]), .C0(n1511_adj_2196[30]), 
          .D0(GND_net), .A1(n38306), .B1(n1412_adj_2194[31]), .C1(n1511_adj_2196[31]), 
          .D1(GND_net), .CIN(n30840), .S0(n1610_adj_2199[30]), .S1(n1610_adj_2199[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_13.INIT0 = 16'h0fff;
    defparam rem_10_add_1043_13.INIT1 = 16'h0fff;
    defparam rem_10_add_1043_13.INJECT1_0 = "NO";
    defparam rem_10_add_1043_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1043_11 (.A0(n1412_adj_2194[28]), .B0(n1511_adj_2196[28]), 
          .C0(GND_net), .D0(n38306), .A1(n38306), .B1(n1412_adj_2194[29]), 
          .C1(n1511_adj_2196[29]), .D1(GND_net), .CIN(n30839), .COUT(n30840), 
          .S0(n1610_adj_2199[28]), .S1(n1610_adj_2199[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_11.INIT0 = 16'hcfc0;
    defparam rem_10_add_1043_11.INIT1 = 16'h0fff;
    defparam rem_10_add_1043_11.INJECT1_0 = "NO";
    defparam rem_10_add_1043_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1043_9 (.A0(n38306), .B0(n1412_adj_2194[26]), .C0(n1511_adj_2196[26]), 
          .D0(GND_net), .A1(n38306), .B1(n1412_adj_2194[27]), .C1(n1511_adj_2196[27]), 
          .D1(GND_net), .CIN(n30838), .COUT(n30839), .S0(n1610_adj_2199[26]), 
          .S1(n1610_adj_2199[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_9.INIT0 = 16'hf000;
    defparam rem_10_add_1043_9.INIT1 = 16'hf000;
    defparam rem_10_add_1043_9.INJECT1_0 = "NO";
    defparam rem_10_add_1043_9.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i20_3_lut_3_lut (.A(pwm_cnt[12]), .B(duty0[12]), 
         .C(n18_adj_1876), .Z(n20_adj_1345)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 rem_10_i1721_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[25]), 
         .D(n2540_adj_1888), .Z(n2639_adj_1388)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1721_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_54_i17_2_lut_rep_376 (.A(pwm_cnt[8]), .B(duty0[8]), 
         .Z(n38381)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i17_2_lut_rep_376.init = 16'h6666;
    CCU2C rem_10_add_1579_3 (.A0(n13616), .B0(n28208), .C0(n2303_adj_2197[13]), 
          .D0(n587), .A1(n13616), .B1(n28208), .C1(n2303_adj_2197[14]), 
          .D1(n2254_adj_1889), .CIN(n31252), .COUT(n31253), .S0(n2402_adj_2198[13]), 
          .S1(n2402_adj_2198[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1579_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1579_3.INJECT1_0 = "NO";
    defparam rem_10_add_1579_3.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_54_i8_3_lut_3_lut (.A(pwm_cnt[8]), .B(duty0[8]), 
         .C(duty0[4]), .Z(n8_adj_1892)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_54_i19_2_lut_rep_377 (.A(pwm_cnt[9]), .B(duty0[9]), 
         .Z(n38382)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i19_2_lut_rep_377.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_54_i16_3_lut_3_lut (.A(pwm_cnt[9]), .B(duty0[9]), 
         .C(n8_adj_1892), .Z(n16_adj_652)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i16_3_lut_3_lut.init = 16'hd4d4;
    CCU2C rem_10_add_1043_7 (.A0(n38306), .B0(n1412_adj_2194[24]), .C0(n1511_adj_2196[24]), 
          .D0(GND_net), .A1(n1412_adj_2194[25]), .B1(n1511_adj_2196[25]), 
          .C1(GND_net), .D1(n38306), .CIN(n30837), .COUT(n30838), .S0(n1610_adj_2199[24]), 
          .S1(n1610_adj_2199[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_7.INIT0 = 16'hf000;
    defparam rem_10_add_1043_7.INIT1 = 16'h303f;
    defparam rem_10_add_1043_7.INJECT1_0 = "NO";
    defparam rem_10_add_1043_7.INJECT1_1 = "NO";
    CCU2C rem_10_add_1579_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n54), .D1(n2[12]), 
          .COUT(n31252), .S1(n2402_adj_2198[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1579_1.INIT0 = 16'h0000;
    defparam rem_10_add_1579_1.INIT1 = 16'habef;
    defparam rem_10_add_1579_1.INJECT1_0 = "NO";
    defparam rem_10_add_1579_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1043_5 (.A0(n1412_adj_2194[22]), .B0(n1511_adj_2196[22]), 
          .C0(n38306), .D0(GND_net), .A1(n38306), .B1(n1412_adj_2194[23]), 
          .C1(n1511_adj_2196[23]), .D1(GND_net), .CIN(n30836), .COUT(n30837), 
          .S0(n1610_adj_2199[22]), .S1(n1610_adj_2199[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_5.INIT0 = 16'h330f;
    defparam rem_10_add_1043_5.INIT1 = 16'hf000;
    defparam rem_10_add_1043_5.INJECT1_0 = "NO";
    defparam rem_10_add_1043_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1043_3 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n38307), .B1(n1511_adj_2196[21]), .C1(n2[19]), .D1(GND_net), 
          .CIN(n30835), .COUT(n30836), .S0(n1610_adj_2199[20]), .S1(n1610_adj_2199[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_3.INIT0 = 16'h2000;
    defparam rem_10_add_1043_3.INIT1 = 16'hcca0;
    defparam rem_10_add_1043_3.INJECT1_0 = "NO";
    defparam rem_10_add_1043_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1043_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n2[19]), 
          .COUT(n30835));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1043_1.INIT0 = 16'h000F;
    defparam rem_10_add_1043_1.INIT1 = 16'hdfff;
    defparam rem_10_add_1043_1.INJECT1_0 = "NO";
    defparam rem_10_add_1043_1.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i9_2_lut_rep_378 (.A(pwm_cnt[4]), .B(duty1[4]), 
         .Z(n38383)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i9_2_lut_rep_378.init = 16'h6666;
    CCU2C rem_10_add_1110_15 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2199[31]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30834), .S0(n1709[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_15.INIT0 = 16'h0f1f;
    defparam rem_10_add_1110_15.INIT1 = 16'h0000;
    defparam rem_10_add_1110_15.INJECT1_0 = "NO";
    defparam rem_10_add_1110_15.INJECT1_1 = "NO";
    LUT4 i31959_3_lut_4_lut (.A(pwm_cnt[4]), .B(duty1[4]), .C(n38387), 
         .D(n38388), .Z(n36795)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i31959_3_lut_4_lut.init = 16'h0009;
    LUT4 pwm_cnt_14__I_0_53_i21_2_lut_rep_379 (.A(pwm_cnt[10]), .B(duty1[10]), 
         .Z(n38384)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i21_2_lut_rep_379.init = 16'h6666;
    CCU2C rem_10_add_1646_21 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[30]), 
          .D0(n38268), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[31]), 
          .D1(n2336_adj_1900), .CIN(n31250), .S0(n2501_adj_2200[30]), 
          .S1(n2501_adj_2200[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_21.INJECT1_0 = "NO";
    defparam rem_10_add_1646_21.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i23_2_lut_rep_380 (.A(pwm_cnt[11]), .B(duty1[11]), 
         .Z(n38385)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i23_2_lut_rep_380.init = 16'h6666;
    LUT4 i31968_2_lut_3_lut_4_lut (.A(pwm_cnt[11]), .B(duty1[11]), .C(duty1[10]), 
         .D(pwm_cnt[10]), .Z(n36804)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i31968_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 pwm_cnt_14__I_0_53_i18_3_lut_3_lut (.A(pwm_cnt[11]), .B(duty1[11]), 
         .C(duty1[10]), .Z(n18_adj_1903)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i18_3_lut_3_lut.init = 16'hd4d4;
    CCU2C rem_10_add_1110_13 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2199[29]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2199[30]), 
          .D1(GND_net), .CIN(n30833), .COUT(n30834), .S0(n1709[29]), 
          .S1(n1709[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1110_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1110_13.INJECT1_0 = "NO";
    defparam rem_10_add_1110_13.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i25_2_lut_rep_381 (.A(pwm_cnt[12]), .B(duty1[12]), 
         .Z(n38386)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i25_2_lut_rep_381.init = 16'h6666;
    CCU2C rem_10_add_1646_19 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[28]), 
          .D0(n2339_adj_1904), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[29]), 
          .D1(n2338_adj_1905), .CIN(n31249), .COUT(n31250), .S0(n2501_adj_2200[28]), 
          .S1(n2501_adj_2200[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_19.INJECT1_0 = "NO";
    defparam rem_10_add_1646_19.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i20_3_lut_3_lut (.A(pwm_cnt[12]), .B(duty1[12]), 
         .C(n18_adj_1903), .Z(n20_adj_1349)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i20_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1646_3 (.A0(n13555), .B0(n28297), .C0(n2402_adj_2195[12]), 
          .D0(n339_adj_1752), .A1(n13555), .B1(n28297), .C1(n2402_adj_2195[13]), 
          .D1(n2354_adj_1910), .CIN(n30700), .COUT(n30701), .S0(n2501_adj_2190[12]), 
          .S1(n2501_adj_2190[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1646_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1646_3.INJECT1_0 = "NO";
    defparam div_9_add_1646_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1110_11 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2199[27]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2199[28]), 
          .D1(n38306), .CIN(n30832), .COUT(n30833), .S0(n1709[27]), 
          .S1(n1709[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_11.INIT0 = 16'hf1e0;
    defparam rem_10_add_1110_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1110_11.INJECT1_0 = "NO";
    defparam rem_10_add_1110_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1110_9 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2199[25]), 
          .D0(n38306), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2199[26]), 
          .D1(GND_net), .CIN(n30831), .COUT(n30832), .S0(n1709[25]), 
          .S1(n1709[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1110_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1110_9.INJECT1_0 = "NO";
    defparam rem_10_add_1110_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1110_7 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2199[23]), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2199[24]), 
          .D1(GND_net), .CIN(n30830), .COUT(n30831), .S0(n1709[23]), 
          .S1(n1709[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_7.INIT0 = 16'hf1e0;
    defparam rem_10_add_1110_7.INIT1 = 16'h0e1f;
    defparam rem_10_add_1110_7.INJECT1_0 = "NO";
    defparam rem_10_add_1110_7.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i17_2_lut_rep_382 (.A(pwm_cnt[8]), .B(duty1[8]), 
         .Z(n38387)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i17_2_lut_rep_382.init = 16'h6666;
    CCU2C div_9_add_976_3 (.A0(n12154), .B0(n5), .C0(n35[19]), .D0(n1412[22]), 
          .A1(n12154), .B1(n5), .C1(n35[19]), .D1(n1412[23]), .CIN(n30612), 
          .COUT(n30613), .S0(n1511_adj_2191[22]), .S1(n1511_adj_2191[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_976_3.INIT0 = 16'h4040;
    defparam div_9_add_976_3.INIT1 = 16'hffff;
    defparam div_9_add_976_3.INJECT1_0 = "NO";
    defparam div_9_add_976_3.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i8_3_lut_3_lut (.A(pwm_cnt[8]), .B(duty1[8]), 
         .C(duty1[4]), .Z(n8_adj_1911)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i8_3_lut_3_lut.init = 16'hd4d4;
    CCU2C div_9_add_1646_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n35[11]), .D1(duty0_14__N_426[9]), 
          .COUT(n30700), .S1(n2501_adj_2190[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1646_1.INIT0 = 16'h0000;
    defparam div_9_add_1646_1.INIT1 = 16'h04bf;
    defparam div_9_add_1646_1.INJECT1_0 = "NO";
    defparam div_9_add_1646_1.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i19_2_lut_rep_383 (.A(pwm_cnt[9]), .B(duty1[9]), 
         .Z(n38388)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i19_2_lut_rep_383.init = 16'h6666;
    CCU2C rem_10_add_1646_17 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[26]), 
          .D0(n2341_adj_1912), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[27]), 
          .D1(n2340_adj_1913), .CIN(n31248), .COUT(n31249), .S0(n2501_adj_2200[26]), 
          .S1(n2501_adj_2200[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_17.INJECT1_0 = "NO";
    defparam rem_10_add_1646_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_1110_5 (.A0(GND_net), .B0(GND_net), .C0(n1610_adj_2199[21]), 
          .D0(n38306), .A1(GND_net), .B1(GND_net), .C1(n1610_adj_2199[22]), 
          .D1(n38306), .CIN(n30829), .COUT(n30830), .S0(n1709[21]), 
          .S1(n1709[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_5.INIT0 = 16'h0e1f;
    defparam rem_10_add_1110_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1110_5.INJECT1_0 = "NO";
    defparam rem_10_add_1110_5.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_21 (.A0(n13557), .B0(n28269), .C0(n2303[31]), 
          .D0(n2237_adj_1916), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n30699), .S0(n2402_adj_2195[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_21.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_21.INIT1 = 16'h0000;
    defparam div_9_add_1579_21.INJECT1_0 = "NO";
    defparam div_9_add_1579_21.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_19 (.A0(n13557), .B0(n28269), .C0(n2303[29]), 
          .D0(n2239_adj_1917), .A1(n13557), .B1(n28269), .C1(n2303[30]), 
          .D1(n2238_adj_1918), .CIN(n30698), .COUT(n30699), .S0(n2402_adj_2195[29]), 
          .S1(n2402_adj_2195[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_19.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_19.INIT1 = 16'h0e1f;
    defparam div_9_add_1579_19.INJECT1_0 = "NO";
    defparam div_9_add_1579_19.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_53_i16_3_lut_3_lut (.A(pwm_cnt[9]), .B(duty1[9]), 
         .C(n8_adj_1911), .Z(n16_adj_625)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i1_2_lut_4_lut_adj_192 (.A(n3228), .B(n3293[30]), .C(n38185), 
         .D(n3326_adj_1304), .Z(n36016)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_192.init = 16'hffca;
    CCU2C rem_10_add_1110_3 (.A0(n27382), .B0(n3), .C0(n5), .D0(n2[19]), 
          .A1(n38307), .B1(n1610_adj_2199[20]), .C1(n2[19]), .D1(GND_net), 
          .CIN(n30828), .COUT(n30829), .S0(n1709[19]), .S1(n1709[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_3.INIT0 = 16'h2000;
    defparam rem_10_add_1110_3.INIT1 = 16'hcca0;
    defparam rem_10_add_1110_3.INJECT1_0 = "NO";
    defparam rem_10_add_1110_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1110_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n27382), .B1(n3), .C1(n5), .D1(n2[18]), 
          .COUT(n30828));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1110_1.INIT0 = 16'h000F;
    defparam rem_10_add_1110_1.INIT1 = 16'hdfff;
    defparam rem_10_add_1110_1.INJECT1_0 = "NO";
    defparam rem_10_add_1110_1.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i9_2_lut_rep_384 (.A(pwm_cnt[4]), .B(duty2[4]), 
         .Z(n38389)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i9_2_lut_rep_384.init = 16'h6666;
    LUT4 rem_10_i1730_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[16]), 
         .D(n2549_adj_1920), .Z(n2648_adj_1335)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1730_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1579_17 (.A0(n13557), .B0(n28269), .C0(n2303[27]), 
          .D0(n2241_adj_1921), .A1(n13557), .B1(n28269), .C1(n2303[28]), 
          .D1(n2240_adj_1922), .CIN(n30697), .COUT(n30698), .S0(n2402_adj_2195[27]), 
          .S1(n2402_adj_2195[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_17.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_17.INIT1 = 16'h0e1f;
    defparam div_9_add_1579_17.INJECT1_0 = "NO";
    defparam div_9_add_1579_17.INJECT1_1 = "NO";
    LUT4 rem_10_i1736_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[10]), 
         .D(n590), .Z(n2654_adj_1413)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1736_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_1401_25 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30826), 
          .S0(n4540[23]), .S1(n4540[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_25.INIT0 = 16'hfff0;
    defparam add_1401_25.INIT1 = 16'hfff0;
    defparam add_1401_25.INJECT1_0 = "NO";
    defparam add_1401_25.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_15 (.A0(n13557), .B0(n28269), .C0(n2303[25]), 
          .D0(n2243_adj_1924), .A1(n13557), .B1(n28269), .C1(n2303[26]), 
          .D1(n2242_adj_1925), .CIN(n30696), .COUT(n30697), .S0(n2402_adj_2195[25]), 
          .S1(n2402_adj_2195[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_15.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_15.INIT1 = 16'h0e1f;
    defparam div_9_add_1579_15.INJECT1_0 = "NO";
    defparam div_9_add_1579_15.INJECT1_1 = "NO";
    LUT4 i32016_3_lut_4_lut (.A(pwm_cnt[4]), .B(duty2[4]), .C(n38393), 
         .D(n38394), .Z(n36852)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32016_3_lut_4_lut.init = 16'h0009;
    CCU2C add_1401_23 (.A0(n35[19]), .B0(n38307), .C0(GND_net), .D0(VCC_net), 
          .A1(n35[19]), .B1(n38307), .C1(GND_net), .D1(VCC_net), .CIN(n30825), 
          .COUT(n30826), .S0(n4540[21]), .S1(n4540[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_23.INIT0 = 16'hffff;
    defparam add_1401_23.INIT1 = 16'h7777;
    defparam add_1401_23.INJECT1_0 = "NO";
    defparam add_1401_23.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i21_2_lut_rep_385 (.A(pwm_cnt[10]), .B(duty2[10]), 
         .Z(n38390)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i21_2_lut_rep_385.init = 16'h6666;
    LUT4 rem_10_i1727_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[19]), 
         .D(n2546_adj_1927), .Z(n2645_adj_1363)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1727_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1646_15 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[24]), 
          .D0(n2343_adj_1928), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[25]), 
          .D1(n2342_adj_1929), .CIN(n31247), .COUT(n31248), .S0(n2501_adj_2200[24]), 
          .S1(n2501_adj_2200[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_15.INJECT1_0 = "NO";
    defparam rem_10_add_1646_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_1646_13 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[22]), 
          .D0(n2345_adj_1932), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[23]), 
          .D1(n2344_adj_1933), .CIN(n31246), .COUT(n31247), .S0(n2501_adj_2200[22]), 
          .S1(n2501_adj_2200[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_13.INJECT1_0 = "NO";
    defparam rem_10_add_1646_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1646_11 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[20]), 
          .D0(n2347_adj_1936), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[21]), 
          .D1(n2346_adj_1937), .CIN(n31245), .COUT(n31246), .S0(n2501_adj_2200[20]), 
          .S1(n2501_adj_2200[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_11.INJECT1_0 = "NO";
    defparam rem_10_add_1646_11.INJECT1_1 = "NO";
    LUT4 div_9_i2124_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[24]), 
         .D(n3135), .Z(n3234)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1733_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[13]), 
         .D(n2552_adj_1941), .Z(n2651_adj_1369)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1733_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1646_9 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[18]), 
          .D0(n2349_adj_1942), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[19]), 
          .D1(n2348_adj_1943), .CIN(n31244), .COUT(n31245), .S0(n2501_adj_2200[18]), 
          .S1(n2501_adj_2200[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1646_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1646_9.INJECT1_0 = "NO";
    defparam rem_10_add_1646_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1646_7 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[16]), 
          .D0(n2351_adj_1946), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[17]), 
          .D1(n2350_adj_1947), .CIN(n31243), .COUT(n31244), .S0(n2501_adj_2200[16]), 
          .S1(n2501_adj_2200[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1646_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1646_7.INJECT1_0 = "NO";
    defparam rem_10_add_1646_7.INJECT1_1 = "NO";
    LUT4 select_842_Select_8_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[8]), 
         .D(n2983), .Z(duty0_14__N_410[8])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_8_i4_3_lut_4_lut.init = 16'hff10;
    CCU2C rem_10_add_1646_5 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[14]), 
          .D0(n2353_adj_1950), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[15]), 
          .D1(n2352_adj_1951), .CIN(n31242), .COUT(n31243), .S0(n2501_adj_2200[14]), 
          .S1(n2501_adj_2200[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1646_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1646_5.INJECT1_0 = "NO";
    defparam rem_10_add_1646_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1646_3 (.A0(n13546), .B0(n28022), .C0(n2402_adj_2198[12]), 
          .D0(n588), .A1(n13546), .B1(n28022), .C1(n2402_adj_2198[13]), 
          .D1(n2354_adj_1954), .CIN(n31241), .COUT(n31242), .S0(n2501_adj_2200[12]), 
          .S1(n2501_adj_2200[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1646_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1646_3.INJECT1_0 = "NO";
    defparam rem_10_add_1646_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1646_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[11]), .D1(duty0_14__N_426[9]), 
          .COUT(n31241), .S1(n2501_adj_2200[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1646_1.INIT0 = 16'h0000;
    defparam rem_10_add_1646_1.INIT1 = 16'h04bf;
    defparam rem_10_add_1646_1.INJECT1_0 = "NO";
    defparam rem_10_add_1646_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1713_23 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[31]), 
          .D0(n2435_adj_1958), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31240), .S0(n2600_adj_2188[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_23.INIT1 = 16'h0000;
    defparam rem_10_add_1713_23.INJECT1_0 = "NO";
    defparam rem_10_add_1713_23.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i23_2_lut_rep_386 (.A(pwm_cnt[11]), .B(duty2[11]), 
         .Z(n38391)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i23_2_lut_rep_386.init = 16'h6666;
    CCU2C rem_10_add_1713_21 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[29]), 
          .D0(n38260), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[30]), 
          .D1(n38261), .CIN(n31239), .COUT(n31240), .S0(n2600_adj_2188[29]), 
          .S1(n2600_adj_2188[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_21.INJECT1_0 = "NO";
    defparam rem_10_add_1713_21.INJECT1_1 = "NO";
    LUT4 i32025_2_lut_3_lut_4_lut (.A(pwm_cnt[11]), .B(duty2[11]), .C(duty2[10]), 
         .D(pwm_cnt[10]), .Z(n36861)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32025_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 pwm_cnt_14__I_0_52_i18_3_lut_3_lut (.A(pwm_cnt[11]), .B(duty2[11]), 
         .C(duty2[10]), .Z(n18_adj_1962)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_52_i25_2_lut_rep_387 (.A(pwm_cnt[12]), .B(duty2[12]), 
         .Z(n38392)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i25_2_lut_rep_387.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_52_i20_3_lut_3_lut (.A(pwm_cnt[12]), .B(duty2[12]), 
         .C(n18_adj_1962), .Z(n20_adj_1351)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i20_3_lut_3_lut.init = 16'hd4d4;
    CCU2C rem_10_add_1713_19 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[27]), 
          .D0(n2439_adj_1963), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[28]), 
          .D1(n2438_adj_1964), .CIN(n31238), .COUT(n31239), .S0(n2600_adj_2188[27]), 
          .S1(n2600_adj_2188[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_19.INJECT1_0 = "NO";
    defparam rem_10_add_1713_19.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_52_i17_2_lut_rep_388 (.A(pwm_cnt[8]), .B(duty2[8]), 
         .Z(n38393)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i17_2_lut_rep_388.init = 16'h6666;
    LUT4 div_9_i2133_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[15]), 
         .D(n3144), .Z(n3243)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2133_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1713_17 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[25]), 
          .D0(n2441_adj_1966), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[26]), 
          .D1(n2440), .CIN(n31237), .COUT(n31238), .S0(n2600_adj_2188[25]), 
          .S1(n2600_adj_2188[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_17.INJECT1_0 = "NO";
    defparam rem_10_add_1713_17.INJECT1_1 = "NO";
    LUT4 div_9_i2123_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[25]), 
         .D(n3134), .Z(n3233_adj_522)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2136_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[12]), 
         .D(n3147), .Z(n3246_adj_548)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2136_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1713_15 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[23]), 
          .D0(n2443_adj_1968), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[24]), 
          .D1(n2442_adj_1969), .CIN(n31236), .COUT(n31237), .S0(n2600_adj_2188[23]), 
          .S1(n2600_adj_2188[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_15.INJECT1_0 = "NO";
    defparam rem_10_add_1713_15.INJECT1_1 = "NO";
    LUT4 rem_10_i1715_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[31]), 
         .D(n2534_adj_1972), .Z(n2633_adj_1348)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1715_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1713_13 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[21]), 
          .D0(n2445_adj_1973), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[22]), 
          .D1(n2444_adj_1974), .CIN(n31235), .COUT(n31236), .S0(n2600_adj_2188[21]), 
          .S1(n2600_adj_2188[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_13.INJECT1_0 = "NO";
    defparam rem_10_add_1713_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1713_11 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[19]), 
          .D0(n2447_adj_1977), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[20]), 
          .D1(n2446_adj_1978), .CIN(n31234), .COUT(n31235), .S0(n2600_adj_2188[19]), 
          .S1(n2600_adj_2188[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_11.INJECT1_0 = "NO";
    defparam rem_10_add_1713_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1713_9 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[17]), 
          .D0(n2449_adj_1980), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[18]), 
          .D1(n2448_adj_1981), .CIN(n31233), .COUT(n31234), .S0(n2600_adj_2188[17]), 
          .S1(n2600_adj_2188[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1713_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1713_9.INJECT1_0 = "NO";
    defparam rem_10_add_1713_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1713_7 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[15]), 
          .D0(n2451_adj_1984), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[16]), 
          .D1(n2450_adj_1985), .CIN(n31232), .COUT(n31233), .S0(n2600_adj_2188[15]), 
          .S1(n2600_adj_2188[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1713_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1713_7.INJECT1_0 = "NO";
    defparam rem_10_add_1713_7.INJECT1_1 = "NO";
    LUT4 div_9_i2134_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[14]), 
         .D(n3145), .Z(n3244)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2134_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2135_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[13]), 
         .D(n3146), .Z(n3245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2135_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1713_5 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[13]), 
          .D0(n2453_adj_1987), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[14]), 
          .D1(n2452_adj_1988), .CIN(n31231), .COUT(n31232), .S0(n2600_adj_2188[13]), 
          .S1(n2600_adj_2188[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1713_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1713_5.INJECT1_0 = "NO";
    defparam rem_10_add_1713_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1713_3 (.A0(n13599), .B0(n28096), .C0(n2501_adj_2200[11]), 
          .D0(n589), .A1(n13599), .B1(n28096), .C1(n2501_adj_2200[12]), 
          .D1(n2454_adj_1990), .CIN(n31230), .COUT(n31231), .S0(n2600_adj_2188[11]), 
          .S1(n2600_adj_2188[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1713_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1713_3.INJECT1_0 = "NO";
    defparam rem_10_add_1713_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1720_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[26]), 
         .D(n2539_adj_1993), .Z(n2638_adj_1428)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1720_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1713_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[10]), .D1(duty0_14__N_426[8]), 
          .COUT(n31230), .S1(n2600_adj_2188[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1713_1.INIT0 = 16'h0000;
    defparam rem_10_add_1713_1.INIT1 = 16'h04bf;
    defparam rem_10_add_1713_1.INJECT1_0 = "NO";
    defparam rem_10_add_1713_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_23 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[30]), 
          .D0(n2535_adj_1994), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[31]), 
          .D1(n2534_adj_1972), .CIN(n31228), .S0(n2699_adj_2180[30]), 
          .S1(n2699_adj_2180[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_23.INJECT1_0 = "NO";
    defparam rem_10_add_1780_23.INJECT1_1 = "NO";
    LUT4 rem_10_i2069_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[12]), 
         .D(n3048_adj_1692), .Z(n3147_adj_1996)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2069_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_193 (.A(n34666), .B(n34856), .C(n3250), .D(n27858), 
         .Z(n28434)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_193.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_194 (.A(n3247_adj_599), .B(n3248_adj_618), .C(n3249_adj_622), 
         .Z(n34666)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_194.init = 16'h8080;
    LUT4 pwm_cnt_14__I_0_52_i8_3_lut_3_lut (.A(pwm_cnt[8]), .B(duty2[8]), 
         .C(duty2[4]), .Z(n8_adj_1997)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 div_9_i2126_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[22]), 
         .D(n3137), .Z(n3236)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1726_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[20]), 
         .D(n2545_adj_1998), .Z(n2644_adj_1415)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1726_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1717_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[29]), 
         .D(n2536_adj_1999), .Z(n2635_adj_1146)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1717_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1716_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[30]), 
         .D(n2535_adj_1994), .Z(n2634_adj_1377)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1716_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1722_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[24]), 
         .D(n38256), .Z(n2640_adj_1434)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1722_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_52_i19_2_lut_rep_389 (.A(pwm_cnt[9]), .B(duty2[9]), 
         .Z(n38394)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i19_2_lut_rep_389.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_52_i16_3_lut_3_lut (.A(pwm_cnt[9]), .B(duty2[9]), 
         .C(n8_adj_1997), .Z(n16_adj_607)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i16_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_51_i9_2_lut_rep_390 (.A(pwm_cnt[4]), .B(duty3[4]), 
         .Z(n38395)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i9_2_lut_rep_390.init = 16'h6666;
    CCU2C rem_10_add_1780_21 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[28]), 
          .D0(n2537_adj_1498), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[29]), 
          .D1(n2536_adj_1999), .CIN(n31227), .COUT(n31228), .S0(n2699_adj_2180[28]), 
          .S1(n2699_adj_2180[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_21.INJECT1_0 = "NO";
    defparam rem_10_add_1780_21.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_19 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[26]), 
          .D0(n2539_adj_1993), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[27]), 
          .D1(n2538_adj_2000), .CIN(n31226), .COUT(n31227), .S0(n2699_adj_2180[26]), 
          .S1(n2699_adj_2180[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_19.INJECT1_0 = "NO";
    defparam rem_10_add_1780_19.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_17 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[24]), 
          .D0(n38256), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[25]), 
          .D1(n2540_adj_1888), .CIN(n31225), .COUT(n31226), .S0(n2699_adj_2180[24]), 
          .S1(n2699_adj_2180[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_17.INJECT1_0 = "NO";
    defparam rem_10_add_1780_17.INJECT1_1 = "NO";
    CCU2C div_9_add_976_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n27382), .B1(n3), .C1(n5), .D1(n35[19]), .COUT(n30612), 
          .S1(n1511_adj_2191[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_976_1.INIT0 = 16'h0000;
    defparam div_9_add_976_1.INIT1 = 16'hdfff;
    defparam div_9_add_976_1.INJECT1_0 = "NO";
    defparam div_9_add_976_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_15 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[22]), 
          .D0(n2543_adj_2001), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[23]), 
          .D1(n2542_adj_2002), .CIN(n31224), .COUT(n31225), .S0(n2699_adj_2180[22]), 
          .S1(n2699_adj_2180[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_15.INJECT1_0 = "NO";
    defparam rem_10_add_1780_15.INJECT1_1 = "NO";
    LUT4 i32073_3_lut_4_lut (.A(pwm_cnt[4]), .B(duty3[4]), .C(n38399), 
         .D(n38400), .Z(n36909)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32073_3_lut_4_lut.init = 16'h0009;
    LUT4 pwm_cnt_14__I_0_51_i21_2_lut_rep_391 (.A(pwm_cnt[10]), .B(duty3[10]), 
         .Z(n38396)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i21_2_lut_rep_391.init = 16'h6666;
    CCU2C rem_10_add_1780_13 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[20]), 
          .D0(n2545_adj_1998), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[21]), 
          .D1(n2544_adj_2003), .CIN(n31223), .COUT(n31224), .S0(n2699_adj_2180[20]), 
          .S1(n2699_adj_2180[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_13.INJECT1_0 = "NO";
    defparam rem_10_add_1780_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_11 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[18]), 
          .D0(n2547_adj_2004), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[19]), 
          .D1(n2546_adj_1927), .CIN(n31222), .COUT(n31223), .S0(n2699_adj_2180[18]), 
          .S1(n2699_adj_2180[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_11.INJECT1_0 = "NO";
    defparam rem_10_add_1780_11.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_51_i23_2_lut_rep_392 (.A(pwm_cnt[11]), .B(duty3[11]), 
         .Z(n38397)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i23_2_lut_rep_392.init = 16'h6666;
    CCU2C rem_10_add_1780_9 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[16]), 
          .D0(n2549_adj_1920), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[17]), 
          .D1(n2548_adj_2005), .CIN(n31221), .COUT(n31222), .S0(n2699_adj_2180[16]), 
          .S1(n2699_adj_2180[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1780_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1780_9.INJECT1_0 = "NO";
    defparam rem_10_add_1780_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_7 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[14]), 
          .D0(n2551_adj_2006), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[15]), 
          .D1(n2550_adj_2007), .CIN(n31220), .COUT(n31221), .S0(n2699_adj_2180[14]), 
          .S1(n2699_adj_2180[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1780_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1780_7.INJECT1_0 = "NO";
    defparam rem_10_add_1780_7.INJECT1_1 = "NO";
    LUT4 div_9_i2120_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[28]), 
         .D(n3131_adj_1727), .Z(n3230)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2120_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1780_5 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[12]), 
          .D0(n2553_adj_2008), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[13]), 
          .D1(n2552_adj_1941), .CIN(n31219), .COUT(n31220), .S0(n2699_adj_2180[12]), 
          .S1(n2699_adj_2180[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1780_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1780_5.INJECT1_0 = "NO";
    defparam rem_10_add_1780_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1780_3 (.A0(n13601), .B0(n28082), .C0(n2600_adj_2188[10]), 
          .D0(n590), .A1(n13601), .B1(n28082), .C1(n2600_adj_2188[11]), 
          .D1(n2554_adj_2009), .CIN(n31218), .COUT(n31219), .S0(n2699_adj_2180[10]), 
          .S1(n2699_adj_2180[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1780_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1780_3.INJECT1_0 = "NO";
    defparam rem_10_add_1780_3.INJECT1_1 = "NO";
    LUT4 i32082_2_lut_3_lut_4_lut (.A(pwm_cnt[11]), .B(duty3[11]), .C(duty3[10]), 
         .D(pwm_cnt[10]), .Z(n36918)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32082_2_lut_3_lut_4_lut.init = 16'h9009;
    LUT4 rem_10_i2070_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[11]), 
         .D(n3049_adj_1694), .Z(n3148_adj_2011)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2070_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1780_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[9]), .D1(duty0_14__N_426[7]), 
          .COUT(n31218), .S1(n2699_adj_2180[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1780_1.INIT0 = 16'h0000;
    defparam rem_10_add_1780_1.INIT1 = 16'h04bf;
    defparam rem_10_add_1780_1.INJECT1_0 = "NO";
    defparam rem_10_add_1780_1.INJECT1_1 = "NO";
    LUT4 pwm_cnt_14__I_0_51_i18_3_lut_3_lut (.A(pwm_cnt[11]), .B(duty3[11]), 
         .C(duty3[10]), .Z(n18_adj_2012)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i18_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_51_i25_2_lut_rep_393 (.A(pwm_cnt[12]), .B(duty3[12]), 
         .Z(n38398)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i25_2_lut_rep_393.init = 16'h6666;
    LUT4 i23909_3_lut (.A(n597), .B(n3253_adj_1776), .C(n3254_adj_597), 
         .Z(n27858)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23909_3_lut.init = 16'hecec;
    LUT4 pwm_cnt_14__I_0_51_i20_3_lut_3_lut (.A(pwm_cnt[12]), .B(duty3[12]), 
         .C(n18_adj_2012), .Z(n20_adj_1374)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i20_3_lut_3_lut.init = 16'hd4d4;
    LUT4 rem_10_i1729_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[17]), 
         .D(n2548_adj_2005), .Z(n2647_adj_1400)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1729_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_51_i17_2_lut_rep_394 (.A(pwm_cnt[8]), .B(duty3[8]), 
         .Z(n38399)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i17_2_lut_rep_394.init = 16'h6666;
    LUT4 rem_10_i1734_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[12]), 
         .D(n2553_adj_2008), .Z(n2652_adj_1365)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1734_3_lut_4_lut.init = 16'hf1e0;
    LUT4 pwm_cnt_14__I_0_51_i8_3_lut_3_lut (.A(pwm_cnt[8]), .B(duty3[8]), 
         .C(duty3[4]), .Z(n8_adj_2013)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i8_3_lut_3_lut.init = 16'hd4d4;
    LUT4 pwm_cnt_14__I_0_51_i19_2_lut_rep_395 (.A(pwm_cnt[9]), .B(duty3[9]), 
         .Z(n38400)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i19_2_lut_rep_395.init = 16'h6666;
    LUT4 pwm_cnt_14__I_0_51_i16_3_lut_3_lut (.A(pwm_cnt[9]), .B(duty3[9]), 
         .C(n8_adj_2013), .Z(n16_adj_589)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i16_3_lut_3_lut.init = 16'hd4d4;
    CCU2C rem_10_add_1847_25 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[31]), 
          .D0(n2633_adj_1348), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31217), .S0(n2798_adj_2165[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_25.INIT1 = 16'h0000;
    defparam rem_10_add_1847_25.INJECT1_0 = "NO";
    defparam rem_10_add_1847_25.INJECT1_1 = "NO";
    LUT4 div_9_i2122_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[26]), 
         .D(n3133_adj_2014), .Z(n3232)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2122_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_add_1579_13 (.A0(n13557), .B0(n28269), .C0(n2303[23]), 
          .D0(n2245_adj_2015), .A1(n13557), .B1(n28269), .C1(n2303[24]), 
          .D1(n2244_adj_2016), .CIN(n30695), .COUT(n30696), .S0(n2402_adj_2195[23]), 
          .S1(n2402_adj_2195[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_13.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_13.INIT1 = 16'h0e1f;
    defparam div_9_add_1579_13.INJECT1_0 = "NO";
    defparam div_9_add_1579_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1732_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[14]), 
         .D(n2551_adj_2006), .Z(n2650_adj_1356)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1732_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1731_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[15]), 
         .D(n2550_adj_2007), .Z(n2649_adj_1340)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1731_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1719_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[27]), 
         .D(n2538_adj_2000), .Z(n2637_adj_1202)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1719_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2130_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[18]), 
         .D(n3141), .Z(n3240)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2130_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1735_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[11]), 
         .D(n2554_adj_2009), .Z(n2653_adj_1214)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1735_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1724_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[22]), 
         .D(n2543_adj_2001), .Z(n2642_adj_1367)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1724_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_1401_21 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n30824), 
          .COUT(n30825), .S0(n4540[19]), .S1(n4540[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_21.INIT0 = 16'h1111;
    defparam add_1401_21.INIT1 = 16'h1111;
    defparam add_1401_21.INJECT1_0 = "NO";
    defparam add_1401_21.INJECT1_1 = "NO";
    LUT4 rem_10_i1723_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[23]), 
         .D(n2542_adj_2002), .Z(n2641_adj_1371)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1723_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1728_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[18]), 
         .D(n2547_adj_2004), .Z(n2646_adj_1391)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1728_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_195 (.A(n36396), .B(n36404), .C(duty0_14__N_426[5]), 
         .D(n38321), .Z(n12416)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_adj_195.init = 16'h0080;
    LUT4 rem_10_i1725_3_lut_4_lut (.A(n28082), .B(n13601), .C(n2600_adj_2188[21]), 
         .D(n2544_adj_2003), .Z(n2643_adj_1419)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1725_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_196 (.A(duty0_14__N_426[2]), .B(n3), .C(n60_adj_4), 
         .D(n63_adj_10), .Z(n36396)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_196.init = 16'ha888;
    LUT4 i1_2_lut_4_lut_adj_197 (.A(n2546_adj_1234), .B(n2600_adj_2186[19]), 
         .C(n38253), .D(n2642_adj_1302), .Z(n36220)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_197.init = 16'hffca;
    LUT4 i1_4_lut_adj_198 (.A(n36472), .B(n36402), .C(n12154), .D(n36470), 
         .Z(n36404)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_198.init = 16'hc0c4;
    LUT4 i24382_2_lut_rep_248 (.A(n28331), .B(n13553), .Z(n38253)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24382_2_lut_rep_248.init = 16'heeee;
    LUT4 div_9_i1726_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[20]), 
         .D(n2545_adj_1233), .Z(n2644_adj_1168)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1726_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1113_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[30]), 
         .D(n38294), .Z(n1743_adj_1421)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1113_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_199 (.A(n36462), .B(n5), .C(n75_adj_1), .D(distance[0]), 
         .Z(n36472)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(59[11:23])
    defparam i1_4_lut_adj_199.init = 16'hfffe;
    LUT4 i1_4_lut_adj_200 (.A(duty0_14__N_426[9]), .B(n3), .C(n81_adj_15), 
         .D(n72_adj_13), .Z(n36402)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_200.init = 16'ha888;
    LUT4 i1_4_lut_adj_201 (.A(n35288), .B(n35294), .C(n35284), .D(n35290), 
         .Z(n13620)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_201.init = 16'hfffe;
    LUT4 i1_4_lut_adj_202 (.A(n42), .B(n48), .C(n39), .D(n45), .Z(n36470)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(59[11:23])
    defparam i1_4_lut_adj_202.init = 16'hfffe;
    LUT4 i1_2_lut_adj_203 (.A(n51), .B(n54), .Z(n36462)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(59[11:23])
    defparam i1_2_lut_adj_203.init = 16'heeee;
    LUT4 div_9_i1725_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[21]), 
         .D(n2544_adj_1239), .Z(n2643_adj_1167)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1725_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2125_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[23]), 
         .D(n3136), .Z(n3235)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_204 (.A(n1), .B(n13790), .C(n89[0]), .D(n197[13]), 
         .Z(duty3_14__N_488[13])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_204.init = 16'h2000;
    LUT4 div_9_i2131_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[17]), 
         .D(n3142), .Z(n3241_adj_532)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2131_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1735_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[11]), 
         .D(n2554_adj_1273), .Z(n2653_adj_1185)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1735_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1731_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[15]), 
         .D(n2550_adj_1260), .Z(n2649_adj_1171)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1731_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1736_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[10]), 
         .D(n341), .Z(n2654_adj_1186)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1736_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1847_23 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[29]), 
          .D0(n2635_adj_1146), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[30]), 
          .D1(n2634_adj_1377), .CIN(n31216), .COUT(n31217), .S0(n2798_adj_2165[29]), 
          .S1(n2798_adj_2165[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_23.INJECT1_0 = "NO";
    defparam rem_10_add_1847_23.INJECT1_1 = "NO";
    CCU2C rem_10_add_1847_21 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[27]), 
          .D0(n2637_adj_1202), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[28]), 
          .D1(n38250), .CIN(n31215), .COUT(n31216), .S0(n2798_adj_2165[27]), 
          .S1(n2798_adj_2165[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_21.INJECT1_0 = "NO";
    defparam rem_10_add_1847_21.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_11 (.A0(n13557), .B0(n28269), .C0(n2303[21]), 
          .D0(n2247_adj_2017), .A1(n13557), .B1(n28269), .C1(n2303[22]), 
          .D1(n2246_adj_2018), .CIN(n30694), .COUT(n30695), .S0(n2402_adj_2195[21]), 
          .S1(n2402_adj_2195[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_11.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_11.INIT1 = 16'h0e1f;
    defparam div_9_add_1579_11.INJECT1_0 = "NO";
    defparam div_9_add_1579_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_205 (.A(n3131), .B(n3194_adj_2167[28]), .C(n38189), 
         .D(n3241_adj_685), .Z(n35028)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_205.init = 16'hffca;
    LUT4 div_9_i1728_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[18]), 
         .D(n2547_adj_1249), .Z(n2646_adj_1157)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1728_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1718_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[28]), 
         .D(n2537_adj_1236), .Z(n2636_adj_1154)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1718_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i28720_3_lut (.A(n13790), .B(n89[0]), .C(n1), .Z(n2983)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(80[9] 86[16])
    defparam i28720_3_lut.init = 16'h5454;
    LUT4 div_13_i2418_4_lut (.A(n28303), .B(n4990[0]), .C(n3556), .D(n13607), 
         .Z(n197[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i2418_4_lut.init = 16'hcfca;
    LUT4 div_9_i1720_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[26]), 
         .D(n2539_adj_1235), .Z(n2638_adj_1165)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1720_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1730_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[16]), 
         .D(n2549_adj_1251), .Z(n2648_adj_1170)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1730_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_206 (.A(n3235_adj_539), .B(n3246), .C(n3230_adj_1779), 
         .D(n3241), .Z(n35288)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_206.init = 16'hfffe;
    LUT4 div_9_i1733_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[13]), 
         .D(n2552_adj_1261), .Z(n2651_adj_1172)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1733_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1727_3_lut_rep_247_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[19]), 
         .D(n2546_adj_1234), .Z(n38252)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1727_3_lut_rep_247_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1715_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[31]), 
         .D(n2534_adj_1248), .Z(n2633)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1715_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1717_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[29]), 
         .D(n2536_adj_1237), .Z(n2635_adj_1153)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1717_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1244_17 (.A0(n13631), .B0(n28090), .C0(n1808[31]), 
          .D0(n1742_adj_1640), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n30611), .S0(n1907[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1244_17.INIT1 = 16'h0000;
    defparam rem_10_add_1244_17.INJECT1_0 = "NO";
    defparam rem_10_add_1244_17.INJECT1_1 = "NO";
    LUT4 div_9_i1719_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[27]), 
         .D(n2538_adj_1245), .Z(n2637_adj_1166)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1719_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1847_19 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[25]), 
          .D0(n2639_adj_1388), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[26]), 
          .D1(n2638_adj_1428), .CIN(n31214), .COUT(n31215), .S0(n2798_adj_2165[25]), 
          .S1(n2798_adj_2165[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_19.INJECT1_0 = "NO";
    defparam rem_10_add_1847_19.INJECT1_1 = "NO";
    LUT4 div_9_i2132_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[16]), 
         .D(n38201), .Z(n3242)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2132_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1734_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[12]), 
         .D(n2553_adj_1272), .Z(n2652_adj_1174)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1734_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1723_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[23]), 
         .D(n2542_adj_1241), .Z(n2641_adj_1156)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1723_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1847_17 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[23]), 
          .D0(n2641_adj_1371), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[24]), 
          .D1(n2640_adj_1434), .CIN(n31213), .COUT(n31214), .S0(n2798_adj_2165[23]), 
          .S1(n2798_adj_2165[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_17.INJECT1_0 = "NO";
    defparam rem_10_add_1847_17.INJECT1_1 = "NO";
    LUT4 div_9_i2121_3_lut_4_lut (.A(n28588), .B(n13547), .C(n3194[27]), 
         .D(n3132_adj_1728), .Z(n3231)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2121_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2409_3_lut_4_lut (.A(n28331), .B(n13553), .C(n38307), 
         .D(n4540[9]), .Z(n89[9])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_9_i2409_3_lut_4_lut.init = 16'hfe0e;
    CCU2C rem_10_add_1847_15 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[21]), 
          .D0(n2643_adj_1419), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[22]), 
          .D1(n2642_adj_1367), .CIN(n31212), .COUT(n31213), .S0(n2798_adj_2165[21]), 
          .S1(n2798_adj_2165[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_15.INJECT1_0 = "NO";
    defparam rem_10_add_1847_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_1847_13 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[19]), 
          .D0(n2645_adj_1363), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[20]), 
          .D1(n2644_adj_1415), .CIN(n31211), .COUT(n31212), .S0(n2798_adj_2165[19]), 
          .S1(n2798_adj_2165[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_13.INJECT1_0 = "NO";
    defparam rem_10_add_1847_13.INJECT1_1 = "NO";
    LUT4 div_9_i1724_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[22]), 
         .D(n2543_adj_1247), .Z(n2642_adj_1302)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1724_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1716_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[30]), 
         .D(n2535_adj_1246), .Z(n2634_adj_1163)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1716_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1721_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[25]), 
         .D(n2540_adj_1238), .Z(n2639_adj_1164)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1721_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2418_4_lut (.A(n28160), .B(n4540[0]), .C(n38307), .D(n13556), 
         .Z(n89[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i2418_4_lut.init = 16'hcfca;
    LUT4 i1_4_lut_adj_207 (.A(n38307), .B(n33356), .C(n33490), .D(n36654), 
         .Z(n13790)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam i1_4_lut_adj_207.init = 16'hfefc;
    LUT4 div_9_i1732_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[14]), 
         .D(n2551_adj_1259), .Z(n2650_adj_1173)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1732_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1722_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[24]), 
         .D(n2541_adj_1240), .Z(n2640_adj_1162)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1722_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1729_3_lut_4_lut (.A(n28331), .B(n13553), .C(n2600_adj_2186[17]), 
         .D(n2548_adj_1250), .Z(n2647_adj_1169)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1729_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1847_11 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[17]), 
          .D0(n2647_adj_1400), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[18]), 
          .D1(n2646_adj_1391), .CIN(n31210), .COUT(n31211), .S0(n2798_adj_2165[17]), 
          .S1(n2798_adj_2165[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_11.INJECT1_0 = "NO";
    defparam rem_10_add_1847_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_208 (.A(n2336), .B(n2402[31]), .C(n38258), 
         .D(n2436), .Z(n35538)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_208.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_209 (.A(n2341), .B(n2402[26]), .C(n38258), 
         .D(n2442), .Z(n35540)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_209.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_210 (.A(n2442_adj_1969), .B(n2501_adj_2200[24]), 
         .C(n38257), .D(n2539_adj_1993), .Z(n35088)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_210.init = 16'hffca;
    LUT4 i60_4_lut (.A(n25_adj_2019), .B(n36356), .C(n38177), .D(n28_adj_2020), 
         .Z(n28160)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i60_4_lut.init = 16'hca0a;
    CCU2C rem_10_add_1847_9 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[15]), 
          .D0(n2649_adj_1340), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[16]), 
          .D1(n2648_adj_1335), .CIN(n31209), .COUT(n31210), .S0(n2798_adj_2165[15]), 
          .S1(n2798_adj_2165[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1847_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1847_9.INJECT1_0 = "NO";
    defparam rem_10_add_1847_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1847_7 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[13]), 
          .D0(n2651_adj_1369), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[14]), 
          .D1(n2650_adj_1356), .CIN(n31208), .COUT(n31209), .S0(n2798_adj_2165[13]), 
          .S1(n2798_adj_2165[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1847_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1847_7.INJECT1_0 = "NO";
    defparam rem_10_add_1847_7.INJECT1_1 = "NO";
    LUT4 i24151_2_lut_rep_252 (.A(n28096), .B(n13599), .Z(n38257)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24151_2_lut_rep_252.init = 16'heeee;
    LUT4 rem_10_i1655_3_lut_rep_251_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[24]), 
         .D(n2442_adj_1969), .Z(n38256)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1655_3_lut_rep_251_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_211 (.A(n3153_adj_2021), .B(n3194_adj_2175[6]), 
         .C(n38199), .D(n3251), .Z(n34856)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_211.init = 16'hca00;
    CCU2C rem_10_add_1847_5 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[11]), 
          .D0(n2653_adj_1214), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[12]), 
          .D1(n2652_adj_1365), .CIN(n31207), .COUT(n31208), .S0(n2798_adj_2165[11]), 
          .S1(n2798_adj_2165[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1847_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1847_5.INJECT1_0 = "NO";
    defparam rem_10_add_1847_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_1847_3 (.A0(n13606), .B0(n28432), .C0(n2699_adj_2180[9]), 
          .D0(n591), .A1(n13606), .B1(n28432), .C1(n2699_adj_2180[10]), 
          .D1(n2654_adj_1413), .CIN(n31206), .COUT(n31207), .S0(n2798_adj_2165[9]), 
          .S1(n2798_adj_2165[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1847_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1847_3.INJECT1_0 = "NO";
    defparam rem_10_add_1847_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_212 (.A(n3392[8]), .B(n3392[9]), .C(n3392[7]), .Z(n36356)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_212.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_213 (.A(n1), .B(n13790), .C(n89[0]), .D(n197[0]), 
         .Z(duty3_14__N_488[0])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_213.init = 16'h2000;
    LUT4 rem_10_i1668_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[11]), 
         .D(n589), .Z(n2554_adj_2009)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1668_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1847_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n66_adj_9), .D1(n2[8]), 
          .COUT(n31206), .S1(n2798_adj_2165[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1847_1.INIT0 = 16'h0000;
    defparam rem_10_add_1847_1.INIT1 = 16'habef;
    defparam rem_10_add_1847_1.INJECT1_0 = "NO";
    defparam rem_10_add_1847_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_214 (.A(n3392[6]), .B(n3392[4]), .C(n3392[5]), .D(n3392[3]), 
         .Z(n28_adj_2020)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_214.init = 16'heaaa;
    LUT4 rem_10_i1663_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[16]), 
         .D(n2450_adj_1985), .Z(n2549_adj_1920)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1663_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24550_2_lut_rep_194 (.A(n28224), .B(n13619), .Z(n38199)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24550_2_lut_rep_194.init = 16'heeee;
    LUT4 rem_10_i1652_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[27]), 
         .D(n2439_adj_1963), .Z(n2538_adj_2000)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1652_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1660_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[19]), 
         .D(n2447_adj_1977), .Z(n2546_adj_1927)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1660_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1667_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[12]), 
         .D(n2454_adj_1990), .Z(n2553_adj_2008)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1667_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1657_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[22]), 
         .D(n2444_adj_1974), .Z(n2543_adj_2001)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1657_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_215 (.A(n35886), .B(n35882), .C(n37672), .D(n37669), 
         .Z(n13556)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_215.init = 16'hfffe;
    LUT4 rem_10_i1654_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[25]), 
         .D(n2441_adj_1966), .Z(n2540_adj_1888)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1654_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1666_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[13]), 
         .D(n2453_adj_1987), .Z(n2552_adj_1941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1666_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2121_3_lut_rep_186_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[27]), 
         .D(n3132), .Z(n38191)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2121_3_lut_rep_186_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1648_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[31]), 
         .D(n2435_adj_1958), .Z(n2534_adj_1972)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1648_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_216 (.A(n37), .B(n37666), .C(n35856), .D(n55), 
         .Z(n35886)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_216.init = 16'hfffe;
    LUT4 rem_10_i1650_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[29]), 
         .D(n38260), .Z(n2536_adj_1999)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1650_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1662_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[17]), 
         .D(n2449_adj_1980), .Z(n2548_adj_2005)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1662_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_217 (.A(n43), .B(n35854), .C(n35858), .D(n33), 
         .Z(n35882)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_217.init = 16'hfffe;
    LUT4 rem_10_i2142_3_lut_rep_193_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[6]), 
         .D(n3153_adj_2021), .Z(n38198)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2142_3_lut_rep_193_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_218 (.A(n3232), .B(n3293[26]), .C(n38185), 
         .D(n3329_adj_2023), .Z(n36022)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_218.init = 16'hffca;
    LUT4 rem_10_i1656_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[23]), 
         .D(n2443_adj_1968), .Z(n2542_adj_2002)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1656_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1661_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[18]), 
         .D(n2448_adj_1981), .Z(n2547_adj_2004)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1661_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2119_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[29]), 
         .D(n3130_adj_2025), .Z(n3229)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1651_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[28]), 
         .D(n2438_adj_1964), .Z(n2537_adj_1498)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1651_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1659_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[20]), 
         .D(n2446_adj_1978), .Z(n2545_adj_1998)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1659_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1658_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[21]), 
         .D(n2445_adj_1973), .Z(n2544_adj_2003)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1658_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_219 (.A(n3340_adj_1749), .B(n23_adj_1277), .C(n3392[17]), 
         .D(n38177), .Z(n35856)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_219.init = 16'hfcee;
    CCU2C rem_10_add_1914_25 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[30]), 
          .D0(n2733_adj_884), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[31]), 
          .D1(n2732_adj_648), .CIN(n31190), .S0(n2897_adj_2162[30]), .S1(n2897_adj_2162[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_25.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_25.INJECT1_0 = "NO";
    defparam rem_10_add_1914_25.INJECT1_1 = "NO";
    LUT4 rem_10_i1653_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[26]), 
         .D(n2440), .Z(n2539_adj_1993)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1653_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1649_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[30]), 
         .D(n38261), .Z(n2535_adj_1994)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1649_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1914_23 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[28]), 
          .D0(n2735_adj_814), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[29]), 
          .D1(n38242), .CIN(n31189), .COUT(n31190), .S0(n2897_adj_2162[28]), 
          .S1(n2897_adj_2162[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_23.INJECT1_0 = "NO";
    defparam rem_10_add_1914_23.INJECT1_1 = "NO";
    CCU2C rem_10_add_1914_21 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[26]), 
          .D0(n2737_adj_798), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[27]), 
          .D1(n38244), .CIN(n31188), .COUT(n31189), .S0(n2897_adj_2162[26]), 
          .S1(n2897_adj_2162[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_21.INJECT1_0 = "NO";
    defparam rem_10_add_1914_21.INJECT1_1 = "NO";
    LUT4 rem_10_i1665_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[14]), 
         .D(n2452_adj_1988), .Z(n2551_adj_2006)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1665_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_220 (.A(n36250), .B(n2345_adj_1812), .C(n2337_adj_1706), 
         .D(n2336_adj_1708), .Z(n13555)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_220.init = 16'hfffe;
    LUT4 rem_10_i1664_3_lut_4_lut (.A(n28096), .B(n13599), .C(n2501_adj_2200[15]), 
         .D(n2451_adj_1984), .Z(n2550_adj_2007)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1664_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24490_2_lut_rep_253 (.A(n28442), .B(n13630), .Z(n38258)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24490_2_lut_rep_253.init = 16'heeee;
    LUT4 i1_4_lut_adj_221 (.A(n2341_adj_1744), .B(n36246), .C(n36234), 
         .D(n2339_adj_1739), .Z(n36250)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_221.init = 16'hfffe;
    LUT4 i1_4_lut_adj_222 (.A(n2344_adj_1814), .B(n2338_adj_1741), .C(n2340_adj_1746), 
         .D(n2342_adj_1771), .Z(n36246)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_222.init = 16'hfffe;
    LUT4 i1_4_lut_adj_223 (.A(n38183), .B(n21_adj_1113), .C(n3392[26]), 
         .D(n38177), .Z(n35854)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_223.init = 16'hfcee;
    LUT4 i1_4_lut_adj_224 (.A(n2348_adj_1863), .B(n28237), .C(n2347_adj_1830), 
         .D(n2349_adj_1861), .Z(n28297)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_224.init = 16'h8000;
    LUT4 rem_10_i2132_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[16]), 
         .D(n3143_adj_1297), .Z(n3242_adj_588)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2132_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1586_3_lut_rep_250_4_lut (.A(n28442), .B(n13630), .C(n2402[26]), 
         .D(n2341), .Z(n38255)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1586_3_lut_rep_250_4_lut.init = 16'hf1e0;
    LUT4 i24284_4_lut (.A(n2351_adj_1867), .B(n2350_adj_1869), .C(n27976), 
         .D(n2352_adj_1880), .Z(n28237)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24284_4_lut.init = 16'heccc;
    CCU2C rem_10_add_1914_19 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[24]), 
          .D0(n2739_adj_816), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[25]), 
          .D1(n2738_adj_760), .CIN(n31187), .COUT(n31188), .S0(n2897_adj_2162[24]), 
          .S1(n2897_adj_2162[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_19.INJECT1_0 = "NO";
    defparam rem_10_add_1914_19.INJECT1_1 = "NO";
    CCU2C rem_10_add_1914_17 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[22]), 
          .D0(n2741_adj_780), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[23]), 
          .D1(n2740), .CIN(n31186), .COUT(n31187), .S0(n2897_adj_2162[22]), 
          .S1(n2897_adj_2162[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_17.INJECT1_0 = "NO";
    defparam rem_10_add_1914_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_1914_15 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[20]), 
          .D0(n2743_adj_890), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[21]), 
          .D1(n2742_adj_892), .CIN(n31185), .COUT(n31186), .S0(n2897_adj_2162[20]), 
          .S1(n2897_adj_2162[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_15.INJECT1_0 = "NO";
    defparam rem_10_add_1914_15.INJECT1_1 = "NO";
    LUT4 i24026_3_lut (.A(n339_adj_1752), .B(n2353_adj_1878), .C(n2354_adj_1910), 
         .Z(n27976)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24026_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_225 (.A(n3228_adj_582), .B(n35286), .C(n35264), 
         .D(n3243_adj_580), .Z(n35294)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_225.init = 16'hfffe;
    LUT4 div_13_i1592_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[20]), 
         .D(n2347), .Z(n2446)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1592_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1914_13 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[18]), 
          .D0(n2745), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[19]), 
          .D1(n2744_adj_822), .CIN(n31184), .COUT(n31185), .S0(n2897_adj_2162[18]), 
          .S1(n2897_adj_2162[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_13.INJECT1_0 = "NO";
    defparam rem_10_add_1914_13.INJECT1_1 = "NO";
    LUT4 rem_10_i2122_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[26]), 
         .D(n3133_adj_2028), .Z(n3232_adj_1767)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2122_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1596_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[16]), 
         .D(n2351), .Z(n2450)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1596_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1582_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[30]), 
         .D(n2337), .Z(n2436)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1582_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1594_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[18]), 
         .D(n2349), .Z(n2448)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1594_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1595_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[17]), 
         .D(n2350), .Z(n2449)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1595_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_226 (.A(n3329_adj_2023), .B(n63_adj_1305), .C(n3392[28]), 
         .D(n38177), .Z(n35858)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_226.init = 16'hfcee;
    CCU2C rem_10_add_1914_11 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[16]), 
          .D0(n2747_adj_824), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[17]), 
          .D1(n2746_adj_818), .CIN(n31183), .COUT(n31184), .S0(n2897_adj_2162[16]), 
          .S1(n2897_adj_2162[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_11.INJECT1_0 = "NO";
    defparam rem_10_add_1914_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1914_9 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[14]), 
          .D0(n2749_adj_941), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[15]), 
          .D1(n2748_adj_911), .CIN(n31182), .COUT(n31183), .S0(n2897_adj_2162[14]), 
          .S1(n2897_adj_2162[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1914_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1914_9.INJECT1_0 = "NO";
    defparam rem_10_add_1914_9.INJECT1_1 = "NO";
    LUT4 div_13_i1597_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[15]), 
         .D(n2352), .Z(n2451)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1597_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1914_7 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[12]), 
          .D0(n2751_adj_950), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[13]), 
          .D1(n2750_adj_943), .CIN(n31181), .COUT(n31182), .S0(n2897_adj_2162[12]), 
          .S1(n2897_adj_2162[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1914_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1914_7.INJECT1_0 = "NO";
    defparam rem_10_add_1914_7.INJECT1_1 = "NO";
    CCU2C rem_10_add_1914_5 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[10]), 
          .D0(n2753_adj_774), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[11]), 
          .D1(n38246), .CIN(n31180), .COUT(n31181), .S0(n2897_adj_2162[10]), 
          .S1(n2897_adj_2162[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1914_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1914_5.INJECT1_0 = "NO";
    defparam rem_10_add_1914_5.INJECT1_1 = "NO";
    LUT4 div_13_i1590_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[22]), 
         .D(n2345), .Z(n2444)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1590_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1914_3 (.A0(n13626), .B0(n28373), .C0(n2798_adj_2165[8]), 
          .D0(n592), .A1(n13626), .B1(n28373), .C1(n2798_adj_2165[9]), 
          .D1(n2754_adj_945), .CIN(n31179), .COUT(n31180), .S0(n2897_adj_2162[8]), 
          .S1(n2897_adj_2162[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1914_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1914_3.INJECT1_0 = "NO";
    defparam rem_10_add_1914_3.INJECT1_1 = "NO";
    CCU2C rem_10_add_1914_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[7]), .D1(duty0_14__N_426[5]), 
          .COUT(n31179), .S1(n2897_adj_2162[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1914_1.INIT0 = 16'h0000;
    defparam rem_10_add_1914_1.INIT1 = 16'h04bf;
    defparam rem_10_add_1914_1.INJECT1_0 = "NO";
    defparam rem_10_add_1914_1.INJECT1_1 = "NO";
    LUT4 div_13_i1588_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[24]), 
         .D(n38262), .Z(n2442)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1588_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1981_27 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[31]), 
          .D0(n38229), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n31178), .S0(n2996_adj_2193[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_27.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_27.INIT1 = 16'h0000;
    defparam rem_10_add_1981_27.INJECT1_0 = "NO";
    defparam rem_10_add_1981_27.INJECT1_1 = "NO";
    CCU2C rem_10_add_1981_25 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[29]), 
          .D0(n2833), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[30]), 
          .D1(n2832_adj_534), .CIN(n31177), .COUT(n31178), .S0(n2996_adj_2193[29]), 
          .S1(n2996_adj_2193[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_25.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_25.INJECT1_0 = "NO";
    defparam rem_10_add_1981_25.INJECT1_1 = "NO";
    CCU2C rem_10_add_1981_23 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[27]), 
          .D0(n2835), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[28]), 
          .D1(n2834), .CIN(n31176), .COUT(n31177), .S0(n2996_adj_2193[27]), 
          .S1(n2996_adj_2193[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_23.INJECT1_0 = "NO";
    defparam rem_10_add_1981_23.INJECT1_1 = "NO";
    CCU2C rem_10_add_1981_21 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[25]), 
          .D0(n38235), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[26]), 
          .D1(n2836), .CIN(n31175), .COUT(n31176), .S0(n2996_adj_2193[25]), 
          .S1(n2996_adj_2193[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_21.INJECT1_0 = "NO";
    defparam rem_10_add_1981_21.INJECT1_1 = "NO";
    CCU2C rem_10_add_1981_19 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[23]), 
          .D0(n2839), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[24]), 
          .D1(n2838_adj_525), .CIN(n31174), .COUT(n31175), .S0(n2996_adj_2193[23]), 
          .S1(n2996_adj_2193[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_19.INJECT1_0 = "NO";
    defparam rem_10_add_1981_19.INJECT1_1 = "NO";
    LUT4 div_13_i1583_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[29]), 
         .D(n2338), .Z(n2437)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1583_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2124_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[24]), 
         .D(n38206), .Z(n3234_adj_630)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2124_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22729_2_lut_4_lut (.A(n1), .B(n13790), .C(n89[0]), .D(n197[14]), 
         .Z(duty3_14__N_488[14])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i22729_2_lut_4_lut.init = 16'h2000;
    LUT4 i22783_2_lut_4_lut (.A(n1), .B(n13790), .C(n89[0]), .D(n197[7]), 
         .Z(duty3_14__N_488[7])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i22783_2_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_adj_227 (.A(n1), .B(n13790), .C(n89[0]), .D(n197[5]), 
         .Z(duty3_14__N_488[5])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_4_lut_adj_227.init = 16'h2000;
    LUT4 div_13_i1585_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[27]), 
         .D(n2340), .Z(n2439)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1585_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22994_2_lut_4_lut (.A(n1), .B(n13790), .C(n89[0]), .D(n197[2]), 
         .Z(duty3_14__N_488[2])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i22994_2_lut_4_lut.init = 16'h2000;
    CCU2C rem_10_add_1981_17 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[21]), 
          .D0(n2841), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[22]), 
          .D1(n38238), .CIN(n31173), .COUT(n31174), .S0(n2996_adj_2193[21]), 
          .S1(n2996_adj_2193[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_17.INJECT1_0 = "NO";
    defparam rem_10_add_1981_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_1981_15 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[19]), 
          .D0(n2843), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[20]), 
          .D1(n2842), .CIN(n31172), .COUT(n31173), .S0(n2996_adj_2193[19]), 
          .S1(n2996_adj_2193[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_15.INJECT1_0 = "NO";
    defparam rem_10_add_1981_15.INJECT1_1 = "NO";
    LUT4 i23997_2_lut_4_lut (.A(n1), .B(n13790), .C(n89[0]), .D(n197[1]), 
         .Z(duty3_14__N_488[1])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i23997_2_lut_4_lut.init = 16'h2000;
    LUT4 rem_10_i2127_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[21]), 
         .D(n3138_adj_2031), .Z(n3237_adj_542)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2127_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1591_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[21]), 
         .D(n2346), .Z(n2445)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1591_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1581_3_lut_rep_249_4_lut (.A(n28442), .B(n13630), .C(n2402[31]), 
         .D(n2336), .Z(n38254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1581_3_lut_rep_249_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_12_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[12]), .Z(duty1_14__N_458[12])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_12_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 select_844_Select_11_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[11]), .Z(duty1_14__N_458[11])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_11_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 div_13_i1600_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[12]), 
         .D(n339), .Z(n2454)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1600_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1981_13 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[17]), 
          .D0(n2845), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[18]), 
          .D1(n2844), .CIN(n31171), .COUT(n31172), .S0(n2996_adj_2193[17]), 
          .S1(n2996_adj_2193[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_13.INJECT1_0 = "NO";
    defparam rem_10_add_1981_13.INJECT1_1 = "NO";
    LUT4 div_13_i1599_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[13]), 
         .D(n2354), .Z(n2453)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1599_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1587_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[25]), 
         .D(n2342), .Z(n2441)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1587_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1593_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[19]), 
         .D(n2348), .Z(n2447)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1593_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1598_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[14]), 
         .D(n2353), .Z(n2452)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1598_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_10_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[10]), .Z(duty1_14__N_458[10])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_10_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 div_13_i1589_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[23]), 
         .D(n2344), .Z(n2443)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1589_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_9_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[9]), .Z(duty1_14__N_458[9])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_9_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 select_844_Select_6_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[6]), .Z(duty1_14__N_458[6])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_6_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 div_13_i1584_3_lut_4_lut (.A(n28442), .B(n13630), .C(n2402[28]), 
         .D(n2339), .Z(n2438)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1584_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_844_Select_4_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[4]), .Z(duty1_14__N_458[4])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_4_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 div_13_i2407_3_lut_4_lut (.A(n28442), .B(n13630), .C(n3556), 
         .D(n4990[11]), .Z(n197[11])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2407_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i24370_2_lut_rep_254 (.A(n28319), .B(n13554), .Z(n38259)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24370_2_lut_rep_254.init = 16'heeee;
    LUT4 div_9_i1648_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[31]), 
         .D(n2435), .Z(n2534_adj_1248)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1648_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1981_11 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[15]), 
          .D0(n2847), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[16]), 
          .D1(n2846), .CIN(n31170), .COUT(n31171), .S0(n2996_adj_2193[15]), 
          .S1(n2996_adj_2193[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_11.INJECT1_0 = "NO";
    defparam rem_10_add_1981_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_228 (.A(n35790), .B(n35820), .C(n3350_adj_2032), 
         .D(n28172), .Z(n28512)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_228.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_229 (.A(n3348_adj_2033), .B(n3347_adj_1112), .C(n3349_adj_2034), 
         .Z(n35790)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_229.init = 16'h8080;
    CCU2C rem_10_add_1981_9 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[13]), 
          .D0(n2849), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[14]), 
          .D1(n2848_adj_570), .CIN(n31169), .COUT(n31170), .S0(n2996_adj_2193[13]), 
          .S1(n2996_adj_2193[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_1981_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_1981_9.INJECT1_0 = "NO";
    defparam rem_10_add_1981_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_1981_7 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[11]), 
          .D0(n2851), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[12]), 
          .D1(n2850), .CIN(n31168), .COUT(n31169), .S0(n2996_adj_2193[11]), 
          .S1(n2996_adj_2193[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_1981_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_1981_7.INJECT1_0 = "NO";
    defparam rem_10_add_1981_7.INJECT1_1 = "NO";
    LUT4 rem_10_i2118_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[30]), 
         .D(n3129_adj_2036), .Z(n3228_adj_582)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1650_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[29]), 
         .D(n2437_adj_1310), .Z(n2536_adj_1237)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1650_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1659_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[20]), 
         .D(n2446_adj_1313), .Z(n2545_adj_1233)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1659_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1668_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[11]), 
         .D(n340_adj_1326), .Z(n2554_adj_1273)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1668_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_230 (.A(n3352), .B(n3252), .C(n3293[6]), .D(n38185), 
         .Z(n35820)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_230.init = 16'ha088;
    LUT4 rem_10_i2129_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[19]), 
         .D(n3140_adj_2038), .Z(n3239_adj_624)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2129_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1658_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[21]), 
         .D(n2445_adj_1311), .Z(n2544_adj_1239)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1658_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n4559_bdd_4_lut (.A(n38272), .B(n38279), .C(n38284), .D(n38285), 
         .Z(n37596)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n4559_bdd_4_lut.init = 16'hfffe;
    LUT4 div_9_i1664_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[15]), 
         .D(n2451_adj_1323), .Z(n2550_adj_1260)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1664_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_231 (.A(n3230_adj_1779), .B(n3293_adj_2161[28]), 
         .C(n38188), .D(n3340), .Z(n34816)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_231.init = 16'hffca;
    LUT4 div_9_i1660_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[19]), 
         .D(n2447_adj_1320), .Z(n2546_adj_1234)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1660_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24220_3_lut (.A(n349_adj_1742), .B(n3353_adj_1636), .C(n3354_adj_1637), 
         .Z(n28172)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24220_3_lut.init = 16'hecec;
    CCU2C rem_10_add_1981_5 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[9]), 
          .D0(n2853), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[10]), 
          .D1(n38237), .CIN(n31167), .COUT(n31168), .S0(n2996_adj_2193[9]), 
          .S1(n2996_adj_2193[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_1981_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_1981_5.INJECT1_0 = "NO";
    defparam rem_10_add_1981_5.INJECT1_1 = "NO";
    LUT4 rem_10_i2134_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[14]), 
         .D(n3145_adj_2040), .Z(n3244_adj_551)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2134_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1666_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[13]), 
         .D(n2453_adj_1327), .Z(n2552_adj_1261)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1666_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1651_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[28]), 
         .D(n2438_adj_1312), .Z(n2537_adj_1236)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1651_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_232 (.A(n36032), .B(n36036), .C(n36026), .D(n36030), 
         .Z(n13602)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_232.init = 16'hfffe;
    LUT4 div_9_i1661_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[18]), 
         .D(n2448_adj_1321), .Z(n2547_adj_1249)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1661_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_233 (.A(n3336_adj_808), .B(n36016), .C(n36022), 
         .D(n3341_adj_1114), .Z(n36032)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_233.init = 16'hfffe;
    CCU2C rem_10_add_1981_3 (.A0(n13598), .B0(n28307), .C0(n2897_adj_2162[7]), 
          .D0(n593), .A1(n13598), .B1(n28307), .C1(n2897_adj_2162[8]), 
          .D1(n2854), .CIN(n31166), .COUT(n31167), .S0(n2996_adj_2193[7]), 
          .S1(n2996_adj_2193[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_1981_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_1981_3.INJECT1_0 = "NO";
    defparam rem_10_add_1981_3.INJECT1_1 = "NO";
    LUT4 rem_10_i2117_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[31]), 
         .D(n3128_adj_2042), .Z(n3227_adj_584)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2117_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1663_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[16]), 
         .D(n2450_adj_1324), .Z(n2549_adj_1251)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1663_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_234 (.A(n3334_adj_1714), .B(n34510), .C(n3343_adj_1525), 
         .D(n3335_adj_1716), .Z(n36036)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_234.init = 16'hfffe;
    LUT4 i24632_2_lut_rep_180 (.A(n28492), .B(n13629), .Z(n38185)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24632_2_lut_rep_180.init = 16'heeee;
    LUT4 i1_4_lut_adj_235 (.A(n3344_adj_2043), .B(n3330_adj_812), .C(n3345_adj_1715), 
         .D(n3328_adj_2044), .Z(n36026)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_235.init = 16'hfffe;
    LUT4 i1_4_lut_adj_236 (.A(n3337_adj_1526), .B(n3338_adj_2045), .C(n3339_adj_875), 
         .D(n3340_adj_1749), .Z(n36030)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_236.init = 16'hfffe;
    LUT4 div_9_i1667_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[12]), 
         .D(n2454_adj_1328), .Z(n2553_adj_1272)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1667_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_237 (.A(n35568), .B(n35566), .C(n2138_adj_1786), 
         .D(n2140_adj_1790), .Z(n13597)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_237.init = 16'hfffe;
    LUT4 rem_10_i2120_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[28]), 
         .D(n3131_adj_2047), .Z(n3230_adj_1779)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2408_3_lut_rep_162_4_lut (.A(n28319), .B(n13554), .C(n38307), 
         .D(n4540[10]), .Z(n38167)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_9_i2408_3_lut_rep_162_4_lut.init = 16'hfe0e;
    LUT4 i1_4_lut_adj_238 (.A(n2139_adj_1785), .B(n2143_adj_1793), .C(n2145_adj_1797), 
         .D(n2144_adj_1798), .Z(n35568)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_238.init = 16'hfffe;
    CCU2C rem_10_add_1981_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[6]), .D1(duty0_14__N_426[4]), 
          .COUT(n31166), .S1(n2996_adj_2193[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1981_1.INIT0 = 16'h0000;
    defparam rem_10_add_1981_1.INIT1 = 16'h04bf;
    defparam rem_10_add_1981_1.INJECT1_0 = "NO";
    defparam rem_10_add_1981_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_239 (.A(n3332_adj_1527), .B(n3342_adj_1713), .C(n3346_adj_1276), 
         .D(n3333_adj_2048), .Z(n34510)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_239.init = 16'hfffe;
    CCU2C rem_10_add_2048_27 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[30]), 
          .D0(n2931_adj_535), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[31]), 
          .D1(n2930), .CIN(n31164), .S0(n3095_adj_2184[30]), .S1(n3095_adj_2184[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_27.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_27.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_27.INJECT1_0 = "NO";
    defparam rem_10_add_2048_27.INJECT1_1 = "NO";
    CCU2C rem_10_add_2048_25 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[28]), 
          .D0(n38220), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[29]), 
          .D1(n2932), .CIN(n31163), .COUT(n31164), .S0(n3095_adj_2184[28]), 
          .S1(n3095_adj_2184[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_25.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_25.INJECT1_0 = "NO";
    defparam rem_10_add_2048_25.INJECT1_1 = "NO";
    LUT4 div_9_i1652_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[27]), 
         .D(n2439_adj_1317), .Z(n2538_adj_1245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1652_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1656_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[23]), 
         .D(n2443_adj_1319), .Z(n2542_adj_1241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1656_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_240 (.A(n2141_adj_1789), .B(n2146_adj_1804), .C(n2142_adj_1794), 
         .Z(n35566)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_3_lut_adj_240.init = 16'hfefe;
    LUT4 div_9_i1653_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[26]), 
         .D(n38265), .Z(n2539_adj_1235)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1653_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2048_23 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[26]), 
          .D0(n2935), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[27]), 
          .D1(n2934), .CIN(n31162), .COUT(n31163), .S0(n3095_adj_2184[26]), 
          .S1(n3095_adj_2184[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_23.INJECT1_0 = "NO";
    defparam rem_10_add_2048_23.INJECT1_1 = "NO";
    LUT4 div_9_i1662_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[17]), 
         .D(n2449_adj_1322), .Z(n2548_adj_1250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1662_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2048_21 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[24]), 
          .D0(n2937_adj_526), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[25]), 
          .D1(n2936), .CIN(n31161), .COUT(n31162), .S0(n3095_adj_2184[24]), 
          .S1(n3095_adj_2184[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_21.INJECT1_0 = "NO";
    defparam rem_10_add_2048_21.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_241 (.A(n2147_adj_1803), .B(n28158), .C(n2148_adj_1808), 
         .D(n2149_adj_1807), .Z(n28387)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_241.init = 16'h8000;
    CCU2C rem_10_add_2048_19 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[22]), 
          .D0(n2939), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[23]), 
          .D1(n2938), .CIN(n31160), .COUT(n31161), .S0(n3095_adj_2184[22]), 
          .S1(n3095_adj_2184[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_19.INJECT1_0 = "NO";
    defparam rem_10_add_2048_19.INJECT1_1 = "NO";
    CCU2C rem_10_add_2048_17 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[20]), 
          .D0(n38225), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[21]), 
          .D1(n2940), .CIN(n31159), .COUT(n31160), .S0(n3095_adj_2184[20]), 
          .S1(n3095_adj_2184[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_17.INJECT1_0 = "NO";
    defparam rem_10_add_2048_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_2048_15 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[18]), 
          .D0(n2943), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[19]), 
          .D1(n2942), .CIN(n31158), .COUT(n31159), .S0(n3095_adj_2184[18]), 
          .S1(n3095_adj_2184[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_15.INJECT1_0 = "NO";
    defparam rem_10_add_2048_15.INJECT1_1 = "NO";
    LUT4 div_9_i1657_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[22]), 
         .D(n2444_adj_1604), .Z(n2543_adj_1247)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1657_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24206_4_lut (.A(n2151_adj_1815), .B(n2150_adj_1816), .C(n27882), 
         .D(n2152_adj_1820), .Z(n28158)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24206_4_lut.init = 16'heccc;
    LUT4 div_9_i1649_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[30]), 
         .D(n2436_adj_1318), .Z(n2535_adj_1246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1649_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23933_3_lut (.A(n586), .B(n2153_adj_1819), .C(n2154_adj_1823), 
         .Z(n27882)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23933_3_lut.init = 16'hecec;
    LUT4 div_9_i1654_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[25]), 
         .D(n38266), .Z(n2540_adj_1238)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1654_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1655_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[24]), 
         .D(n2442_adj_1601), .Z(n2541_adj_1240)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1655_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2048_13 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[16]), 
          .D0(n2945), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[17]), 
          .D1(n2944), .CIN(n31157), .COUT(n31158), .S0(n3095_adj_2184[16]), 
          .S1(n3095_adj_2184[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_13.INJECT1_0 = "NO";
    defparam rem_10_add_2048_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_2048_11 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[14]), 
          .D0(n2947_adj_571), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[15]), 
          .D1(n2946), .CIN(n31156), .COUT(n31157), .S0(n3095_adj_2184[14]), 
          .S1(n3095_adj_2184[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_11.INJECT1_0 = "NO";
    defparam rem_10_add_2048_11.INJECT1_1 = "NO";
    LUT4 div_9_i1665_3_lut_4_lut (.A(n28319), .B(n13554), .C(n2501_adj_2190[14]), 
         .D(n2452_adj_1325), .Z(n2551_adj_1259)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1665_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2133_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[15]), 
         .D(n3144_adj_2067), .Z(n3243_adj_580)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2133_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_242 (.A(n2338_adj_1905), .B(n2402_adj_2198[29]), 
         .C(n38264), .D(n2445_adj_1973), .Z(n35590)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_242.init = 16'hffca;
    CCU2C rem_10_add_2048_9 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[12]), 
          .D0(n2949), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[13]), 
          .D1(n2948), .CIN(n31155), .COUT(n31156), .S0(n3095_adj_2184[12]), 
          .S1(n3095_adj_2184[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_2048_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_2048_9.INJECT1_0 = "NO";
    defparam rem_10_add_2048_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_243 (.A(n38268), .B(n2402_adj_2198[30]), .C(n38264), 
         .D(n2438_adj_1964), .Z(n35588)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_243.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_244 (.A(n2244), .B(n2303_adj_2171[24]), .C(n38263), 
         .D(n2345), .Z(n35608)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_244.init = 16'hffca;
    LUT4 rem_10_i2123_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[25]), 
         .D(n3134_adj_2070), .Z(n3233)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2123_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_245 (.A(n35584), .B(n35582), .C(n2241_adj_1836), 
         .D(n2245_adj_1844), .Z(n13616)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_245.init = 16'hfffe;
    LUT4 div_9_i2185_3_lut_rep_176_4_lut (.A(n28492), .B(n13629), .C(n3293[30]), 
         .D(n3228), .Z(n38181)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2185_3_lut_rep_176_4_lut.init = 16'hf1e0;
    LUT4 i24484_2_lut_rep_258 (.A(n28430), .B(n13633), .Z(n38263)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24484_2_lut_rep_258.init = 16'heeee;
    CCU2C rem_10_add_2048_7 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[10]), 
          .D0(n2951), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[11]), 
          .D1(n2950), .CIN(n31154), .COUT(n31155), .S0(n3095_adj_2184[10]), 
          .S1(n3095_adj_2184[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_2048_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_2048_7.INJECT1_0 = "NO";
    defparam rem_10_add_2048_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_246 (.A(n2246_adj_1849), .B(n2240_adj_1837), .C(n2243_adj_1840), 
         .D(n2244_adj_1845), .Z(n35584)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_246.init = 16'hfffe;
    LUT4 i1_4_lut_adj_247 (.A(n2238_adj_1833), .B(n2237_adj_1827), .C(n2242_adj_1841), 
         .D(n2239_adj_1832), .Z(n35582)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_247.init = 16'hfffe;
    LUT4 div_9_i2189_3_lut_rep_178_4_lut (.A(n28492), .B(n13629), .C(n3293[26]), 
         .D(n3232), .Z(n38183)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2189_3_lut_rep_178_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_248 (.A(n2247_adj_1848), .B(n28154), .C(n2248_adj_1853), 
         .D(n2249_adj_1852), .Z(n28208)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_248.init = 16'h8000;
    LUT4 i24202_4_lut (.A(n2251_adj_1856), .B(n2250_adj_1857), .C(n27876), 
         .D(n2252_adj_1873), .Z(n28154)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24202_4_lut.init = 16'heccc;
    LUT4 rem_10_i2135_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[13]), 
         .D(n3146_adj_2073), .Z(n3245_adj_642)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2135_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_249 (.A(n35900), .B(n31386), .C(n35902), .D(n35898), 
         .Z(n33356)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_249.init = 16'hfffe;
    LUT4 i23927_3_lut (.A(n587), .B(n2253_adj_1872), .C(n2254_adj_1889), 
         .Z(n27876)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23927_3_lut.init = 16'hecec;
    LUT4 div_13_i1526_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[19]), 
         .D(n2249), .Z(n2348)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1526_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2130_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[18]), 
         .D(n3141_adj_2075), .Z(n3240_adj_561)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2130_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1519_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[26]), 
         .D(n2242), .Z(n2341)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1519_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_1401_19 (.A0(n28287), .B0(n13653), .C0(GND_net), .D0(VCC_net), 
          .A1(GND_net), .B1(n38305), .C1(GND_net), .D1(VCC_net), .CIN(n30823), 
          .COUT(n30824), .S0(n4540[17]), .S1(n4540[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_19.INIT0 = 16'h1111;
    defparam add_1401_19.INIT1 = 16'h1111;
    defparam add_1401_19.INJECT1_0 = "NO";
    defparam add_1401_19.INJECT1_1 = "NO";
    CCU2C rem_10_add_2048_5 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[8]), 
          .D0(n2953), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[9]), 
          .D1(n38224), .CIN(n31153), .COUT(n31154), .S0(n3095_adj_2184[8]), 
          .S1(n3095_adj_2184[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_2048_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_2048_5.INJECT1_0 = "NO";
    defparam rem_10_add_2048_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_2048_3 (.A0(n13592), .B0(n28436), .C0(n2996_adj_2193[6]), 
          .D0(n594), .A1(n13592), .B1(n28436), .C1(n2996_adj_2193[7]), 
          .D1(n2954), .CIN(n31152), .COUT(n31153), .S0(n3095_adj_2184[6]), 
          .S1(n3095_adj_2184[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_2048_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_2048_3.INJECT1_0 = "NO";
    defparam rem_10_add_2048_3.INJECT1_1 = "NO";
    CCU2C add_1401_17 (.A0(n28526), .B0(n13613), .C0(GND_net), .D0(VCC_net), 
          .A1(n28321), .B1(n38289), .C1(GND_net), .D1(VCC_net), .CIN(n30822), 
          .COUT(n30823), .S0(n4540[15]), .S1(n4540[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_17.INIT0 = 16'h1111;
    defparam add_1401_17.INIT1 = 16'h1111;
    defparam add_1401_17.INJECT1_0 = "NO";
    defparam add_1401_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_250 (.A(n35940), .B(n37597), .C(n38418), .D(n35938), 
         .Z(n33490)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam i1_4_lut_adj_250.init = 16'hfffe;
    LUT4 rem_10_i2128_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[20]), 
         .D(n3139_adj_2080), .Z(n3238_adj_639)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2128_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2048_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n75_adj_1), .D1(n2[5]), 
          .COUT(n31152), .S1(n3095_adj_2184[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2048_1.INIT0 = 16'h0000;
    defparam rem_10_add_2048_1.INIT1 = 16'habef;
    defparam rem_10_add_2048_1.INJECT1_0 = "NO";
    defparam rem_10_add_2048_1.INJECT1_1 = "NO";
    CCU2C add_1401_15 (.A0(n28440), .B0(n13590), .C0(GND_net), .D0(VCC_net), 
          .A1(n28263), .B1(n13605), .C1(GND_net), .D1(VCC_net), .CIN(n30821), 
          .COUT(n30822), .S0(n4540[13]), .S1(n4540[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_15.INIT0 = 16'h1111;
    defparam add_1401_15.INIT1 = 16'h1111;
    defparam add_1401_15.INJECT1_0 = "NO";
    defparam add_1401_15.INJECT1_1 = "NO";
    LUT4 div_9_i2206_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[9]), 
         .D(n3249), .Z(n3348_adj_2033)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2206_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1525_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[20]), 
         .D(n2248), .Z(n2347)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1525_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_251 (.A(n38267), .B(n89[7]), .C(n4540[11]), .D(n38307), 
         .Z(n35940)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam i1_4_lut_adj_251.init = 16'hfcee;
    LUT4 rem_10_i2136_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[12]), 
         .D(n3147_adj_1996), .Z(n3246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2136_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_1244_15 (.A0(n13631), .B0(n28090), .C0(n1808[29]), 
          .D0(n1744), .A1(n13631), .B1(n28090), .C1(n1808[30]), .D1(n1743_adj_1643), 
          .CIN(n30610), .COUT(n30611), .S0(n1907[29]), .S1(n1907[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_1244_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_1244_15.INJECT1_0 = "NO";
    defparam rem_10_add_1244_15.INJECT1_1 = "NO";
    LUT4 div_13_i1529_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[16]), 
         .D(n2252), .Z(n2351)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1529_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i26582_4_lut (.A(n38306), .B(n34956), .C(n34958), .D(n1709[31]), 
         .Z(n13631)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i26582_4_lut.init = 16'haaa8;
    LUT4 div_9_i2208_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[7]), 
         .D(n38196), .Z(n3350_adj_2032)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2208_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2115_29 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[31]), 
          .D0(n38210), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n31151), .S0(n3194_adj_2175[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_29.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_29.INIT1 = 16'h0000;
    defparam rem_10_add_2115_29.INJECT1_0 = "NO";
    defparam rem_10_add_2115_29.INJECT1_1 = "NO";
    CCU2C rem_10_add_2115_27 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[29]), 
          .D0(n3031_adj_1629), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[30]), 
          .D1(n3030_adj_1665), .CIN(n31150), .COUT(n31151), .S0(n3194_adj_2175[29]), 
          .S1(n3194_adj_2175[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_27.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_27.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_27.INJECT1_0 = "NO";
    defparam rem_10_add_2115_27.INJECT1_1 = "NO";
    LUT4 div_13_i1527_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[18]), 
         .D(n2250), .Z(n2349)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1527_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_252 (.A(n38247), .B(n89[6]), .C(n4540[8]), .D(n38307), 
         .Z(n35938)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam i1_4_lut_adj_252.init = 16'hfcee;
    LUT4 div_13_i1528_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[17]), 
         .D(n2251), .Z(n2350)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1528_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2115_25 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[27]), 
          .D0(n3033_adj_1670), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[28]), 
          .D1(n3032_adj_1642), .CIN(n31149), .COUT(n31150), .S0(n3194_adj_2175[27]), 
          .S1(n3194_adj_2175[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_25.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_25.INJECT1_0 = "NO";
    defparam rem_10_add_2115_25.INJECT1_1 = "NO";
    CCU2C rem_10_add_2115_23 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[25]), 
          .D0(n3035_adj_1657), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[26]), 
          .D1(n3034_adj_1677), .CIN(n31148), .COUT(n31149), .S0(n3194_adj_2175[25]), 
          .S1(n3194_adj_2175[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_23.INJECT1_0 = "NO";
    defparam rem_10_add_2115_23.INJECT1_1 = "NO";
    LUT4 div_13_i1515_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[30]), 
         .D(n2238), .Z(n2337)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1515_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2115_21 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[23]), 
          .D0(n3037_adj_1667), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[24]), 
          .D1(n3036_adj_1673), .CIN(n31147), .COUT(n31148), .S0(n3194_adj_2175[23]), 
          .S1(n3194_adj_2175[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_21.INJECT1_0 = "NO";
    defparam rem_10_add_2115_21.INJECT1_1 = "NO";
    LUT4 div_13_i1523_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[22]), 
         .D(n2246), .Z(n2345)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1523_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_253 (.A(n35534), .B(n35526), .C(n35532), .D(n2338_adj_1905), 
         .Z(n13546)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_253.init = 16'hfffe;
    CCU2C rem_10_add_2115_19 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[21]), 
          .D0(n3039_adj_1663), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[22]), 
          .D1(n38215), .CIN(n31146), .COUT(n31147), .S0(n3194_adj_2175[21]), 
          .S1(n3194_adj_2175[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_19.INJECT1_0 = "NO";
    defparam rem_10_add_2115_19.INJECT1_1 = "NO";
    CCU2C rem_10_add_2115_17 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[19]), 
          .D0(n3041_adj_1675), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[20]), 
          .D1(n3040_adj_1645), .CIN(n31145), .COUT(n31146), .S0(n3194_adj_2175[19]), 
          .S1(n3194_adj_2175[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_17.INJECT1_0 = "NO";
    defparam rem_10_add_2115_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_2115_15 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[17]), 
          .D0(n3043_adj_1639), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[18]), 
          .D1(n3042_adj_1653), .CIN(n31144), .COUT(n31145), .S0(n3194_adj_2175[17]), 
          .S1(n3194_adj_2175[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_15.INJECT1_0 = "NO";
    defparam rem_10_add_2115_15.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_254 (.A(n2340_adj_1913), .B(n2336_adj_1900), .C(n2343_adj_1928), 
         .D(n2344_adj_1933), .Z(n35534)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_254.init = 16'hfffe;
    LUT4 i1_4_lut_adj_255 (.A(n2339_adj_1904), .B(n2346_adj_1937), .C(n2345_adj_1932), 
         .D(n2342_adj_1929), .Z(n35532)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_255.init = 16'hfffe;
    LUT4 i1_4_lut_adj_256 (.A(n2347_adj_1936), .B(n27996), .C(n2348_adj_1943), 
         .D(n2349_adj_1942), .Z(n28022)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_256.init = 16'h8000;
    LUT4 select_844_Select_3_i3_2_lut_4_lut (.A(n89[0]), .B(n13790), .C(n1), 
         .D(n197[3]), .Z(duty1_14__N_458[3])) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_3_i3_2_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_158 (.A(n89[0]), .B(n13790), .Z(n38163)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam i1_2_lut_rep_158.init = 16'heeee;
    LUT4 i24046_4_lut (.A(n2351_adj_1946), .B(n2350_adj_1947), .C(n27745), 
         .D(n2352_adj_1951), .Z(n27996)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24046_4_lut.init = 16'heccc;
    LUT4 i23799_3_lut (.A(n588), .B(n2353_adj_1950), .C(n2354_adj_1954), 
         .Z(n27745)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23799_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_257 (.A(n36264), .B(n36262), .C(n2240_adj_1922), 
         .D(n2246_adj_2018), .Z(n13557)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_257.init = 16'hfffe;
    LUT4 i1_4_lut_adj_258 (.A(n2241_adj_1921), .B(n2238_adj_1918), .C(n2239_adj_1917), 
         .D(n2242_adj_1925), .Z(n36264)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_258.init = 16'hfffe;
    CCU2C rem_10_add_2115_13 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[15]), 
          .D0(n3045_adj_1633), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[16]), 
          .D1(n3044_adj_1296), .CIN(n31143), .COUT(n31144), .S0(n3194_adj_2175[15]), 
          .S1(n3194_adj_2175[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_13.INJECT1_0 = "NO";
    defparam rem_10_add_2115_13.INJECT1_1 = "NO";
    CCU2C rem_10_add_2115_11 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[13]), 
          .D0(n3047_adj_1690), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[14]), 
          .D1(n3046_adj_1651), .CIN(n31142), .COUT(n31143), .S0(n3194_adj_2175[13]), 
          .S1(n3194_adj_2175[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_11.INJECT1_0 = "NO";
    defparam rem_10_add_2115_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_259 (.A(n2243_adj_1924), .B(n2237_adj_1916), .C(n2244_adj_2016), 
         .D(n2245_adj_2015), .Z(n36262)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_259.init = 16'hfffe;
    LUT4 i1_4_lut_adj_260 (.A(n2247_adj_2017), .B(n28241), .C(n2248_adj_2086), 
         .D(n2249_adj_2087), .Z(n28269)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_260.init = 16'h8000;
    CCU2C rem_10_add_2115_9 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[11]), 
          .D0(n3049_adj_1694), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[12]), 
          .D1(n3048_adj_1692), .CIN(n31141), .COUT(n31142), .S0(n3194_adj_2175[11]), 
          .S1(n3194_adj_2175[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_2115_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_2115_9.INJECT1_0 = "NO";
    defparam rem_10_add_2115_9.INJECT1_1 = "NO";
    LUT4 i24288_4_lut (.A(n2251_adj_2089), .B(n2250_adj_2090), .C(n27982), 
         .D(n2252_adj_2091), .Z(n28241)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24288_4_lut.init = 16'heccc;
    LUT4 i24032_3_lut (.A(n338), .B(n2253_adj_2092), .C(n2254_adj_2093), 
         .Z(n27982)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24032_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_261 (.A(n35606), .B(n2441_adj_1966), .C(n35590), 
         .D(n2443_adj_1968), .Z(n13599)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_261.init = 16'hfffe;
    LUT4 div_9_i2210_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[5]), 
         .D(n3253), .Z(n3352)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2210_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2115_7 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[9]), 
          .D0(n3051_adj_1624), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[10]), 
          .D1(n3050_adj_1700), .CIN(n31140), .COUT(n31141), .S0(n3194_adj_2175[9]), 
          .S1(n3194_adj_2175[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_2115_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_2115_7.INJECT1_0 = "NO";
    defparam rem_10_add_2115_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_262 (.A(n2442_adj_1969), .B(n35602), .C(n35588), 
         .D(n2435_adj_1958), .Z(n35606)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_262.init = 16'hfffe;
    LUT4 i1_4_lut_adj_263 (.A(n2439_adj_1963), .B(n2440), .C(n2446_adj_1978), 
         .D(n2444_adj_1974), .Z(n35602)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_263.init = 16'hfffe;
    LUT4 div_13_i1524_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[21]), 
         .D(n2247), .Z(n2346)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1524_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_264 (.A(n2447_adj_1977), .B(n27988), .C(n2448_adj_1981), 
         .D(n2449_adj_1980), .Z(n28096)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_264.init = 16'h8000;
    LUT4 i24038_4_lut (.A(n2451_adj_1984), .B(n2450_adj_1985), .C(n27735), 
         .D(n2452_adj_1988), .Z(n27988)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24038_4_lut.init = 16'heccc;
    LUT4 i23789_3_lut (.A(n589), .B(n2453_adj_1987), .C(n2454_adj_1990), 
         .Z(n27735)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23789_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_265 (.A(n35096), .B(n35060), .C(n2543_adj_2001), 
         .D(n2540_adj_1888), .Z(n13601)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_265.init = 16'hfffe;
    LUT4 div_13_i1530_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[15]), 
         .D(n2253), .Z(n2352)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1530_3_lut_4_lut.init = 16'hf1e0;
    LUT4 select_842_Select_12_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[12]), .D(n1), .Z(duty0_14__N_410[12])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_12_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 rem_10_i2126_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[22]), 
         .D(n3137_adj_2096), .Z(n3236_adj_568)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2126_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1518_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[27]), 
         .D(n2241), .Z(n2340)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1518_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1514_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[31]), 
         .D(n2237), .Z(n2336)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1514_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_266 (.A(n2546_adj_1927), .B(n35092), .C(n35088), 
         .D(n2545_adj_1998), .Z(n35096)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_266.init = 16'hfffe;
    LUT4 i1_3_lut_adj_267 (.A(n2538_adj_2000), .B(n2535_adj_1994), .C(n2537_adj_1498), 
         .Z(n35060)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_3_lut_adj_267.init = 16'hfefe;
    LUT4 i1_4_lut_adj_268 (.A(n2536_adj_1999), .B(n2544_adj_2003), .C(n2534_adj_1972), 
         .D(n2542_adj_2002), .Z(n35092)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_268.init = 16'hfffe;
    LUT4 rem_10_i2125_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[23]), 
         .D(n3136_adj_2097), .Z(n3235_adj_539)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2125_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_269 (.A(n2547_adj_2004), .B(n27970), .C(n2548_adj_2005), 
         .D(n2549_adj_1920), .Z(n28082)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_269.init = 16'h8000;
    CCU2C rem_10_add_2115_5 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[7]), 
          .D0(n3053_adj_1679), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[8]), 
          .D1(n38216), .CIN(n31139), .COUT(n31140), .S0(n3194_adj_2175[7]), 
          .S1(n3194_adj_2175[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_2115_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_2115_5.INJECT1_0 = "NO";
    defparam rem_10_add_2115_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_2115_3 (.A0(n13628), .B0(n28281), .C0(n3095_adj_2184[5]), 
          .D0(n595), .A1(n13628), .B1(n28281), .C1(n3095_adj_2184[6]), 
          .D1(n3054_adj_1686), .CIN(n31138), .COUT(n31139), .S0(n3194_adj_2175[5]), 
          .S1(n3194_adj_2175[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_2115_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_2115_3.INJECT1_0 = "NO";
    defparam rem_10_add_2115_3.INJECT1_1 = "NO";
    LUT4 i24020_4_lut (.A(n2551_adj_2006), .B(n2550_adj_2007), .C(n27199), 
         .D(n2552_adj_1941), .Z(n27970)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24020_4_lut.init = 16'heccc;
    LUT4 i1_4_lut_adj_270 (.A(n3227_adj_584), .B(n3237_adj_542), .C(n3242_adj_588), 
         .D(n3236_adj_568), .Z(n35284)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_270.init = 16'hfffe;
    LUT4 i23256_3_lut (.A(n590), .B(n2553_adj_2008), .C(n2554_adj_2009), 
         .Z(n27199)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23256_3_lut.init = 16'hecec;
    LUT4 rem_10_i2131_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[17]), 
         .D(n3142_adj_2101), .Z(n3241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2131_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_271 (.A(n38204), .B(n89[2]), .C(n4540[4]), .D(n38307), 
         .Z(n35898)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_271.init = 16'hfcee;
    LUT4 div_13_i1516_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[29]), 
         .D(n2239), .Z(n2338)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1516_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1521_3_lut_rep_257_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[24]), 
         .D(n2244), .Z(n38262)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1521_3_lut_rep_257_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_272 (.A(n35648), .B(n35642), .C(n2642_adj_1367), 
         .D(n2635_adj_1146), .Z(n13606)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_272.init = 16'hfffe;
    LUT4 i1_4_lut_adj_273 (.A(n2633_adj_1348), .B(n35644), .C(n35636), 
         .D(n2646_adj_1391), .Z(n35648)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_273.init = 16'hfffe;
    CCU2C rem_10_add_2115_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[4]), .D1(duty0_14__N_426[2]), 
          .COUT(n31138), .S1(n3194_adj_2175[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2115_1.INIT0 = 16'h0000;
    defparam rem_10_add_2115_1.INIT1 = 16'h04bf;
    defparam rem_10_add_2115_1.INJECT1_0 = "NO";
    defparam rem_10_add_2115_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_274 (.A(n2639_adj_1388), .B(n2638_adj_1428), .C(n2643_adj_1419), 
         .D(n2640_adj_1434), .Z(n35642)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_274.init = 16'hfffe;
    LUT4 i1_4_lut_adj_275 (.A(n2645_adj_1363), .B(n2641_adj_1371), .C(n2634_adj_1377), 
         .D(n2637_adj_1202), .Z(n35644)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_275.init = 16'hfffe;
    LUT4 i1_4_lut_adj_276 (.A(n34804), .B(n5_adj_2103), .C(n13_adj_1564), 
         .D(n27994), .Z(n28303)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_276.init = 16'hc8c0;
    LUT4 select_842_Select_11_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[11]), .D(n1), .Z(duty0_14__N_410[11])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_11_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 div_13_i1532_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[13]), 
         .D(n338_adj_913), .Z(n2354)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1532_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_277 (.A(n38174), .B(n3452_adj_1559), .C(n3392_adj_2177[5]), 
         .D(n38168), .Z(n34804)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_277.init = 16'hc088;
    LUT4 i24044_4_lut (.A(n27749), .B(n3354_adj_1736), .C(n3392_adj_2177[3]), 
         .D(n38168), .Z(n27994)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i24044_4_lut.init = 16'hfaee;
    LUT4 div_13_i1531_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[14]), 
         .D(n2254), .Z(n2353)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1531_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_278 (.A(n2647_adj_1400), .B(n28192), .C(n2648_adj_1335), 
         .D(n2649_adj_1340), .Z(n28432)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_278.init = 16'h8000;
    LUT4 div_13_i1522_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[23]), 
         .D(n2245), .Z(n2344)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1522_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1520_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[25]), 
         .D(n2243), .Z(n2342)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1520_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23803_4_lut (.A(n138), .B(n3454_adj_1548), .C(n38[1]), .D(n3556), 
         .Z(n27749)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i23803_4_lut.init = 16'hc088;
    LUT4 div_13_i1517_3_lut_4_lut (.A(n28430), .B(n13633), .C(n2303_adj_2171[28]), 
         .D(n2240), .Z(n2339)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1517_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24240_4_lut (.A(n2651_adj_1369), .B(n2650_adj_1356), .C(n27923), 
         .D(n2652_adj_1365), .Z(n28192)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24240_4_lut.init = 16'heccc;
    LUT4 div_13_i2406_3_lut_4_lut (.A(n28430), .B(n13633), .C(n3556), 
         .D(n4990[12]), .Z(n197[12])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2406_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i23973_3_lut (.A(n591), .B(n2653_adj_1214), .C(n2654_adj_1413), 
         .Z(n27923)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23973_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_279 (.A(n37517), .B(n35130), .C(n35132), .D(n37506), 
         .Z(n13607)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_279.init = 16'hfffe;
    LUT4 div_9_i2184_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[31]), 
         .D(n3227), .Z(n3326_adj_1304)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_280 (.A(n23_adj_1510), .B(n35102), .C(n35106), .D(n31_adj_1517), 
         .Z(n35130)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_280.init = 16'hfffe;
    LUT4 i1_4_lut_adj_281 (.A(n47), .B(n37488), .C(n35110), .D(n43_adj_1522), 
         .Z(n35132)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_281.init = 16'hfffe;
    LUT4 div_9_i2196_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[19]), 
         .D(n3239), .Z(n3338_adj_2045)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2196_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2143_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[5]), 
         .D(n3154_adj_2106), .Z(n3253_adj_1776)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2143_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2182_29 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[30]), 
          .D0(n3129_adj_2036), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[31]), 
          .D1(n3128_adj_2042), .CIN(n31136), .S0(n3293_adj_2161[30]), 
          .S1(n3293_adj_2161[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_29.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_29.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_29.INJECT1_0 = "NO";
    defparam rem_10_add_2182_29.INJECT1_1 = "NO";
    CCU2C rem_10_add_2182_27 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[28]), 
          .D0(n3131_adj_2047), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[29]), 
          .D1(n3130_adj_2025), .CIN(n31135), .COUT(n31136), .S0(n3293_adj_2161[28]), 
          .S1(n3293_adj_2161[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_27.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_27.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_27.INJECT1_0 = "NO";
    defparam rem_10_add_2182_27.INJECT1_1 = "NO";
    PFUMX i32273 (.BLUT(n37516), .ALUT(n37515), .C0(n38168), .Z(n37517));
    LUT4 select_842_Select_10_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[10]), .D(n1), .Z(duty0_14__N_410[10])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_10_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 select_842_Select_9_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[9]), .D(n1), .Z(duty0_14__N_410[9])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_9_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i24230_2_lut_rep_259 (.A(n28022), .B(n13546), .Z(n38264)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24230_2_lut_rep_259.init = 16'heeee;
    LUT4 i1_4_lut_adj_282 (.A(n35498), .B(n35496), .C(n39_adj_523), .D(n31), 
         .Z(n33697)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_282.init = 16'hfffe;
    LUT4 select_842_Select_6_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[6]), .D(n1), .Z(duty0_14__N_410[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_6_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_283 (.A(n38171), .B(n35494), .C(n35486), .D(n3435), 
         .Z(n35498)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_283.init = 16'hfffe;
    LUT4 select_842_Select_4_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[4]), .D(n1), .Z(duty0_14__N_410[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_4_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_284 (.A(n3446), .B(n3437), .C(n3440), .D(n3436), 
         .Z(n35496)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_284.init = 16'hfffe;
    LUT4 i1_4_lut_adj_285 (.A(n53_adj_1542), .B(n3340_adj_1655), .C(n3392_adj_2177[17]), 
         .D(n38168), .Z(n35102)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_285.init = 16'hfaee;
    LUT4 i1_4_lut_adj_286 (.A(n63_adj_1575), .B(n3344_adj_721), .C(n3392_adj_2177[13]), 
         .D(n38168), .Z(n35106)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_286.init = 16'hfaee;
    LUT4 i1_4_lut_adj_287 (.A(n3434), .B(n3443), .C(n3441), .D(n38169), 
         .Z(n35494)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_287.init = 16'hfffe;
    LUT4 i1_4_lut_adj_288 (.A(n2748), .B(n28289), .C(n2747), .D(n2749), 
         .Z(n28468)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_288.init = 16'h8000;
    LUT4 i24336_4_lut (.A(n2751), .B(n2750), .C(n28040), .D(n2752), 
         .Z(n28289)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24336_4_lut.init = 16'heccc;
    CCU2C rem_10_add_2182_25 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[26]), 
          .D0(n3133_adj_2028), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[27]), 
          .D1(n3132), .CIN(n31134), .COUT(n31135), .S0(n3293_adj_2161[26]), 
          .S1(n3293_adj_2161[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_25.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_25.INJECT1_0 = "NO";
    defparam rem_10_add_2182_25.INJECT1_1 = "NO";
    LUT4 div_9_i2191_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[24]), 
         .D(n3234), .Z(n3333_adj_2048)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_289 (.A(n3329), .B(n49), .C(n3392_adj_2177[28]), 
         .D(n38168), .Z(n35110)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_289.init = 16'hfcee;
    LUT4 i24090_3_lut (.A(n343), .B(n2753), .C(n2754), .Z(n28040)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24090_3_lut.init = 16'hecec;
    LUT4 select_842_Select_3_i3_2_lut_3_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n197[3]), .D(n1), .Z(duty0_14__N_410[3])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(81[11:12])
    defparam select_842_Select_3_i3_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_290 (.A(n35376), .B(n35394), .C(n35392), .D(n2736), 
         .Z(n13622)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_290.init = 16'hfffe;
    LUT4 select_844_Select_1_i4_3_lut_4_lut_4_lut (.A(n89[0]), .B(n13790), 
         .C(n1), .D(n197[1]), .Z(duty1_14__N_458[1])) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A (B+!(C)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(82[11:12])
    defparam select_844_Select_1_i4_3_lut_4_lut_4_lut.init = 16'h3230;
    LUT4 i1_3_lut_4_lut_adj_291 (.A(n38164), .B(n33356), .C(n36350), .D(n1), 
         .Z(n13642)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_291.init = 16'hfeff;
    LUT4 rem_10_i1583_3_lut_rep_255_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[29]), 
         .D(n2338_adj_1905), .Z(n38260)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1583_3_lut_rep_255_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_292 (.A(n2739), .B(n35390), .C(n35384), .D(n2734), 
         .Z(n35394)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_292.init = 16'hfffe;
    LUT4 i1_4_lut_adj_293 (.A(n2744), .B(n2733), .C(n2732), .D(n2737), 
         .Z(n35392)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_293.init = 16'hfffe;
    CCU2C rem_10_add_2182_23 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[24]), 
          .D0(n38206), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[25]), 
          .D1(n3134_adj_2070), .CIN(n31133), .COUT(n31134), .S0(n3293_adj_2161[24]), 
          .S1(n3293_adj_2161[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_23.INJECT1_0 = "NO";
    defparam rem_10_add_2182_23.INJECT1_1 = "NO";
    CCU2C rem_10_add_2182_21 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[22]), 
          .D0(n3137_adj_2096), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[23]), 
          .D1(n3136_adj_2097), .CIN(n31132), .COUT(n31133), .S0(n3293_adj_2161[22]), 
          .S1(n3293_adj_2161[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_21.INJECT1_0 = "NO";
    defparam rem_10_add_2182_21.INJECT1_1 = "NO";
    CCU2C rem_10_add_2182_19 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[20]), 
          .D0(n3139_adj_2080), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[21]), 
          .D1(n3138_adj_2031), .CIN(n31131), .COUT(n31132), .S0(n3293_adj_2161[20]), 
          .S1(n3293_adj_2161[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_19.INJECT1_0 = "NO";
    defparam rem_10_add_2182_19.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_294 (.A(n2743), .B(n2741), .C(n2746), .D(n2742), 
         .Z(n35390)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_294.init = 16'hfffe;
    LUT4 rem_10_i1582_3_lut_rep_256_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[30]), 
         .D(n38268), .Z(n38261)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1582_3_lut_rep_256_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1593_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[19]), 
         .D(n2348_adj_1943), .Z(n2447_adj_1977)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1593_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1596_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[16]), 
         .D(n2351_adj_1946), .Z(n2450_adj_1985)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1596_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_rep_160 (.A(n4540[22]), .B(n4540[21]), .C(n4540[19]), 
         .Z(n38165)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_160.init = 16'hfefe;
    LUT4 i1_2_lut_4_lut_adj_295 (.A(n4540[22]), .B(n4540[21]), .C(n4540[19]), 
         .D(n4540[24]), .Z(n36654)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_295.init = 16'hfffe;
    LUT4 rem_10_i1600_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[12]), 
         .D(n588), .Z(n2454_adj_1990)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1600_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_296 (.A(n2948_adj_1550), .B(n28279), .C(n2947_adj_1620), 
         .D(n2949_adj_1552), .Z(n28506)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_296.init = 16'h8000;
    LUT4 i24326_4_lut (.A(n2951_adj_1514), .B(n2950_adj_1616), .C(n28024), 
         .D(n2952_adj_2110), .Z(n28279)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24326_4_lut.init = 16'heccc;
    LUT4 rem_10_i1585_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[27]), 
         .D(n2340_adj_1913), .Z(n2439_adj_1963)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1585_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24074_3_lut (.A(n345_adj_2111), .B(n2953_adj_1586), .C(n2954_adj_2112), 
         .Z(n28024)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24074_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_297 (.A(n35262), .B(n35252), .C(n2945_adj_1590), 
         .D(n2938_adj_1618), .Z(n13618)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_297.init = 16'hfffe;
    LUT4 i1_4_lut_adj_298 (.A(n35260), .B(n2942_adj_1592), .C(n2930_adj_1583), 
         .D(n2940_adj_1501), .Z(n35262)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_298.init = 16'hfffe;
    CCU2C rem_10_add_2182_17 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[18]), 
          .D0(n3141_adj_2075), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[19]), 
          .D1(n3140_adj_2038), .CIN(n31130), .COUT(n31131), .S0(n3293_adj_2161[18]), 
          .S1(n3293_adj_2161[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_17.INJECT1_0 = "NO";
    defparam rem_10_add_2182_17.INJECT1_1 = "NO";
    CCU2C rem_10_add_2182_15 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[16]), 
          .D0(n3143_adj_1297), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[17]), 
          .D1(n3142_adj_2101), .CIN(n31129), .COUT(n31130), .S0(n3293_adj_2161[16]), 
          .S1(n3293_adj_2161[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_15.INJECT1_0 = "NO";
    defparam rem_10_add_2182_15.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_299 (.A(n2939_adj_1579), .B(n2934_adj_1556), .C(n2937_adj_2113), 
         .D(n2936_adj_1577), .Z(n35252)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_299.init = 16'hfffe;
    LUT4 i1_4_lut_adj_300 (.A(n2935_adj_2114), .B(n35254), .C(n35240), 
         .D(n2933), .Z(n35260)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_300.init = 16'hfffe;
    LUT4 i1_4_lut_adj_301 (.A(n34912), .B(n34904), .C(n3350_adj_1649), 
         .D(n28002), .Z(n28267)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_301.init = 16'ha8a0;
    CCU2C add_1401_13 (.A0(n28297), .B0(n13555), .C0(GND_net), .D0(VCC_net), 
          .A1(n28269), .B1(n13557), .C1(GND_net), .D1(VCC_net), .CIN(n30820), 
          .COUT(n30821), .S0(n4540[11]), .S1(n4540[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_13.INIT0 = 16'h1111;
    defparam add_1401_13.INIT1 = 16'h1111;
    defparam add_1401_13.INJECT1_0 = "NO";
    defparam add_1401_13.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_302 (.A(n3349_adj_1724), .B(n3347_adj_1210), .C(n3348_adj_1757), 
         .Z(n34912)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_302.init = 16'h8080;
    LUT4 i24052_3_lut (.A(n349), .B(n3353_adj_1558), .C(n3354_adj_1736), 
         .Z(n28002)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24052_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_303 (.A(n35334), .B(n35330), .C(n35322), .D(n35324), 
         .Z(n13608)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_303.init = 16'hfffe;
    LUT4 i1_4_lut_adj_304 (.A(n35328), .B(n3342_adj_1516), .C(n3333_adj_1572), 
         .D(n3336_adj_1521), .Z(n35334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_304.init = 16'hfffe;
    LUT4 i1_4_lut_adj_305 (.A(n2931_adj_2115), .B(n2946_adj_2116), .C(n2943_adj_1588), 
         .D(n2944_adj_2117), .Z(n35254)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_305.init = 16'hfffe;
    CCU2C rem_10_add_2182_13 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[14]), 
          .D0(n3145_adj_2040), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[15]), 
          .D1(n3144_adj_2067), .CIN(n31128), .COUT(n31129), .S0(n3293_adj_2161[14]), 
          .S1(n3293_adj_2161[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_13.INJECT1_0 = "NO";
    defparam rem_10_add_2182_13.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_306 (.A(n3338_adj_1307), .B(n35318), .C(n35302), 
         .D(n3327_adj_632), .Z(n35330)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_306.init = 16'hfffe;
    CCU2C rem_10_add_2182_11 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[12]), 
          .D0(n3147_adj_1996), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[13]), 
          .D1(n3146_adj_2073), .CIN(n31127), .COUT(n31128), .S0(n3293_adj_2161[12]), 
          .S1(n3293_adj_2161[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_11.INJECT1_0 = "NO";
    defparam rem_10_add_2182_11.INJECT1_1 = "NO";
    LUT4 rem_10_i2144_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[4]), 
         .D(n596), .Z(n3254_adj_597)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2144_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_307 (.A(n3340_adj_1655), .B(n3335_adj_635), .C(n3332_adj_633), 
         .D(n3334_adj_1561), .Z(n35322)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_307.init = 16'hfffe;
    LUT4 i1_4_lut_adj_308 (.A(n2848_adj_646), .B(n28285), .C(n2847_adj_610), 
         .D(n2849_adj_631), .Z(n28484)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_308.init = 16'h8000;
    LUT4 i24332_4_lut (.A(n2851_adj_647), .B(n2850_adj_636), .C(n28030), 
         .D(n2852), .Z(n28285)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24332_4_lut.init = 16'heccc;
    LUT4 i1_4_lut_adj_309 (.A(n3328_adj_1306), .B(n3346_adj_1509), .C(n3329), 
         .D(n3343_adj_1209), .Z(n35324)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_309.init = 16'hfffe;
    LUT4 i1_4_lut_adj_310 (.A(n3326_adj_1574), .B(n3344_adj_721), .C(n3345_adj_634), 
         .D(n3339_adj_565), .Z(n35328)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_310.init = 16'hfffe;
    LUT4 i24080_3_lut (.A(n344_adj_2118), .B(n2853_adj_591), .C(n2854_adj_601), 
         .Z(n28030)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24080_3_lut.init = 16'hecec;
    LUT4 rem_10_i1590_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[22]), 
         .D(n2345_adj_1932), .Z(n2444_adj_1974)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1590_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2182_9 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[10]), 
          .D0(n3149_adj_2119), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[11]), 
          .D1(n3148_adj_2011), .CIN(n31126), .COUT(n31127), .S0(n3293_adj_2161[10]), 
          .S1(n3293_adj_2161[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_2182_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_2182_9.INJECT1_0 = "NO";
    defparam rem_10_add_2182_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_2182_7 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[8]), 
          .D0(n3151_adj_1294), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[9]), 
          .D1(n3150_adj_2120), .CIN(n31125), .COUT(n31126), .S0(n3293_adj_2161[8]), 
          .S1(n3293_adj_2161[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_2182_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_2182_7.INJECT1_0 = "NO";
    defparam rem_10_add_2182_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_311 (.A(n35468), .B(n35476), .C(n35452), .D(n35462), 
         .Z(n13621)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_311.init = 16'hfffe;
    LUT4 i1_4_lut_adj_312 (.A(n2841_adj_616), .B(n2837), .C(n2835_adj_619), 
         .D(n2832_adj_592), .Z(n35468)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_312.init = 16'hfffe;
    LUT4 i1_4_lut_adj_313 (.A(n2831), .B(n35472), .C(n35466), .D(n2842_adj_620), 
         .Z(n35476)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_313.init = 16'hfffe;
    LUT4 rem_10_i1599_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[13]), 
         .D(n2354_adj_1954), .Z(n2453_adj_1987)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1599_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2141_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[7]), 
         .D(n38205), .Z(n3251)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2141_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_314 (.A(n2836_adj_628), .B(n2834_adj_640), .C(n2846_adj_615), 
         .D(n2843_adj_637), .Z(n35472)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_314.init = 16'hfffe;
    LUT4 rem_10_i1591_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[21]), 
         .D(n2346_adj_1937), .Z(n2445_adj_1973)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1591_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1581_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[31]), 
         .D(n2336_adj_1900), .Z(n2435_adj_1958)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1581_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i8_3_lut (.A(n120), .B(n38[7]), .C(n3556), .Z(n344_adj_2118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i8_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1595_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[17]), 
         .D(n2350_adj_1947), .Z(n2449_adj_1980)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1595_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_315 (.A(n3148_adj_810), .B(n28271), .C(n3147_adj_770), 
         .D(n3149_adj_694), .Z(n28522)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_315.init = 16'h8000;
    LUT4 i24318_4_lut (.A(n3151), .B(n3150_adj_697), .C(n28014), .D(n3152_adj_671), 
         .Z(n28271)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24318_4_lut.init = 16'heccc;
    LUT4 i24064_3_lut (.A(n347_adj_667), .B(n3153_adj_717), .C(n3154_adj_656), 
         .Z(n28014)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24064_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_316 (.A(n35368), .B(n35366), .C(n35348), .D(n3146_adj_768), 
         .Z(n13614)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_316.init = 16'hfffe;
    LUT4 i1_4_lut_adj_317 (.A(n3136_adj_791), .B(n35362), .C(n35342), 
         .D(n3133), .Z(n35368)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_317.init = 16'hfffe;
    LUT4 rem_10_i1584_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[28]), 
         .D(n2339_adj_1904), .Z(n2438_adj_1964)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1584_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2137_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[11]), 
         .D(n3148_adj_2011), .Z(n3247_adj_599)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2137_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_318 (.A(n3128), .B(n35358), .C(n35338), .D(n3135_adj_687), 
         .Z(n35366)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_318.init = 16'hfffe;
    LUT4 i1_4_lut_adj_319 (.A(n3238_adj_639), .B(n3233), .C(n3245_adj_642), 
         .D(n3239_adj_624), .Z(n35290)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_319.init = 16'hfffe;
    LUT4 rem_10_i1586_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[26]), 
         .D(n2341_adj_1912), .Z(n2440)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1586_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_320 (.A(n3134_adj_794), .B(n3144_adj_691), .C(n3141_adj_730), 
         .D(n3140_adj_772), .Z(n35362)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_320.init = 16'hfffe;
    LUT4 i1_4_lut_adj_321 (.A(n3142_adj_684), .B(n3131), .C(n3145_adj_806), 
         .D(n3138_adj_661), .Z(n35358)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_321.init = 16'hfffe;
    LUT4 i1_4_lut_adj_322 (.A(n3048_adj_1404), .B(n28277), .C(n3047_adj_1398), 
         .D(n3049_adj_1483), .Z(n28518)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_322.init = 16'h8000;
    LUT4 i24324_4_lut (.A(n3051_adj_1382), .B(n3050_adj_1181), .C(n28018), 
         .D(n3052_adj_1373), .Z(n28277)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24324_4_lut.init = 16'heccc;
    LUT4 rem_10_i1587_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[25]), 
         .D(n2342_adj_1929), .Z(n2441_adj_1966)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1587_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1594_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[18]), 
         .D(n2349_adj_1942), .Z(n2448_adj_1981)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1594_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24068_3_lut (.A(n346_adj_1140), .B(n3053_adj_1183), .C(n3054_adj_1265), 
         .Z(n28018)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24068_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_323 (.A(n35050), .B(n35000), .C(n34998), .D(n34988), 
         .Z(n13617)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_323.init = 16'hfffe;
    LUT4 i1_4_lut_adj_324 (.A(n3042_adj_1299), .B(n35046), .C(n35042), 
         .D(n3037_adj_1475), .Z(n35050)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_324.init = 16'hfffe;
    CCU2C rem_10_add_2182_5 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[6]), 
          .D0(n3153_adj_2021), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[7]), 
          .D1(n38205), .CIN(n31124), .COUT(n31125), .S0(n3293_adj_2161[6]), 
          .S1(n3293_adj_2161[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_2182_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_2182_5.INJECT1_0 = "NO";
    defparam rem_10_add_2182_5.INJECT1_1 = "NO";
    CCU2C rem_10_add_2182_3 (.A0(n13619), .B0(n28224), .C0(n3194_adj_2175[4]), 
          .D0(n596), .A1(n13619), .B1(n28224), .C1(n3194_adj_2175[5]), 
          .D1(n3154_adj_2106), .CIN(n31123), .COUT(n31124), .S0(n3293_adj_2161[4]), 
          .S1(n3293_adj_2161[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_2182_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_2182_3.INJECT1_0 = "NO";
    defparam rem_10_add_2182_3.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_325 (.A(n3043_adj_1354), .B(n3031), .C(n3036_adj_1176), 
         .D(n3045_adj_1217), .Z(n35000)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_325.init = 16'hfffe;
    LUT4 i1_4_lut_adj_326 (.A(n3032_adj_1417), .B(n3029_adj_1316), .C(n3030), 
         .D(n3039_adj_1358), .Z(n34998)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_326.init = 16'hfffe;
    LUT4 i1_4_lut_adj_327 (.A(n3038_adj_1227), .B(n3033_adj_1055), .C(n3035_adj_1469), 
         .D(n3044_adj_1386), .Z(n35046)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_327.init = 16'hfffe;
    LUT4 rem_10_i2138_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[10]), 
         .D(n3149_adj_2119), .Z(n3248_adj_618)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2138_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n4559_bdd_4_lut_32291 (.A(n4540[13]), .B(n4540[15]), .C(n4540[14]), 
         .D(n4540[16]), .Z(n37595)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n4559_bdd_4_lut_32291.init = 16'hfffe;
    LUT4 n3395_bdd_4_lut (.A(n3328_adj_2044), .B(n3344_adj_2043), .C(n3333_adj_2048), 
         .D(n3338_adj_2045), .Z(n37668)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam n3395_bdd_4_lut.init = 16'hfffe;
    LUT4 select_842_Select_7_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[7]), 
         .D(n2983), .Z(duty0_14__N_410[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_7_i4_3_lut_4_lut.init = 16'hff10;
    LUT4 rem_10_i1589_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[23]), 
         .D(n2344_adj_1933), .Z(n2443_adj_1968)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1589_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1588_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[24]), 
         .D(n2343_adj_1928), .Z(n2442_adj_1969)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1588_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1597_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[15]), 
         .D(n2352_adj_1951), .Z(n2451_adj_1984)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1597_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2204_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[11]), 
         .D(n3247), .Z(n3346_adj_1276)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2204_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_328 (.A(n3248_adj_695), .B(n28261), .C(n3247_adj_811), 
         .D(n3249_adj_698), .Z(n28528)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_328.init = 16'h8000;
    LUT4 i24308_4_lut (.A(n3251_adj_672), .B(n3250_adj_704), .C(n28010), 
         .D(n3252_adj_718), .Z(n28261)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24308_4_lut.init = 16'heccc;
    CCU2C rem_10_add_2182_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n2[3]), .D1(duty0_14__N_426[1]), 
          .COUT(n31123), .S1(n3293_adj_2161[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2182_1.INIT0 = 16'h0000;
    defparam rem_10_add_2182_1.INIT1 = 16'h04bf;
    defparam rem_10_add_2182_1.INJECT1_0 = "NO";
    defparam rem_10_add_2182_1.INJECT1_1 = "NO";
    CCU2C rem_10_add_2249_31 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[31]), 
          .D0(n3227_adj_584), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31122), .S0(n3392_adj_2163[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_31.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_31.INIT1 = 16'h0000;
    defparam rem_10_add_2249_31.INJECT1_0 = "NO";
    defparam rem_10_add_2249_31.INJECT1_1 = "NO";
    LUT4 i24060_3_lut (.A(n348_adj_1735), .B(n3253_adj_657), .C(n3254_adj_668), 
         .Z(n28010)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24060_3_lut.init = 16'hecec;
    LUT4 rem_10_i1592_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[20]), 
         .D(n2347_adj_1936), .Z(n2446_adj_1978)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1592_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_329 (.A(n35036), .B(n35020), .C(n35016), .D(n35018), 
         .Z(n13610)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_329.init = 16'hfffe;
    LUT4 i1_4_lut_adj_330 (.A(n3237_adj_662), .B(n35032), .C(n35028), 
         .D(n3227_adj_726), .Z(n35036)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_330.init = 16'hfffe;
    LUT4 i1_4_lut_adj_331 (.A(n3235_adj_792), .B(n3246_adj_736), .C(n3233_adj_795), 
         .D(n3244_adj_807), .Z(n35020)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_331.init = 16'hfffe;
    CCU2C rem_10_add_2249_29 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[29]), 
          .D0(n3229), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[30]), 
          .D1(n3228_adj_582), .CIN(n31121), .COUT(n31122), .S0(n3392_adj_2163[29]), 
          .S1(n3392_adj_2163[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_29.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_29.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_29.INJECT1_0 = "NO";
    defparam rem_10_add_2249_29.INJECT1_1 = "NO";
    LUT4 rem_10_i1598_3_lut_4_lut (.A(n28022), .B(n13546), .C(n2402_adj_2198[14]), 
         .D(n2353_adj_1950), .Z(n2452_adj_1988)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1598_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2139_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[9]), 
         .D(n3150_adj_2120), .Z(n3249_adj_622)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2139_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i18_3_lut (.A(n90), .B(n38[17]), .C(n3556), .Z(n334_adj_1199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i18_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_332 (.A(n3238_adj_754), .B(n3234_adj_688), .C(n3243_adj_692), 
         .D(n3232_adj_766), .Z(n35016)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_332.init = 16'hfffe;
    LUT4 i1_4_lut_adj_333 (.A(n3236_adj_675), .B(n3229_adj_723), .C(n3242_adj_603), 
         .D(n3231_adj_612), .Z(n35018)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_333.init = 16'hfffe;
    LUT4 i1_4_lut_adj_334 (.A(n3228_adj_682), .B(n3240_adj_564), .C(n3245_adj_720), 
         .D(n3239_adj_773), .Z(n35032)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_334.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_335 (.A(n2341_adj_1744), .B(n2402_adj_2195[26]), 
         .C(n38267), .D(n2442_adj_1601), .Z(n36270)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_335.init = 16'hffca;
    CCU2C rem_10_add_2249_27 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[27]), 
          .D0(n38191), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[28]), 
          .D1(n3230_adj_1779), .CIN(n31120), .COUT(n31121), .S0(n3392_adj_2163[27]), 
          .S1(n3392_adj_2163[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_27.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_27.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_27.INJECT1_0 = "NO";
    defparam rem_10_add_2249_27.INJECT1_1 = "NO";
    CCU2C rem_10_add_2249_25 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[25]), 
          .D0(n3233), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[26]), 
          .D1(n3232_adj_1767), .CIN(n31119), .COUT(n31120), .S0(n3392_adj_2163[25]), 
          .S1(n3392_adj_2163[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_25.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_25.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_25.INJECT1_0 = "NO";
    defparam rem_10_add_2249_25.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_336 (.A(n36650), .B(n38167), .C(n4540[24]), .D(n4540[1]), 
         .Z(n35976)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_336.init = 16'h0100;
    LUT4 rem_10_i2140_3_lut_4_lut (.A(n28224), .B(n13619), .C(n3194_adj_2175[8]), 
         .D(n3151_adj_1294), .Z(n3250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2140_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2202_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[13]), 
         .D(n3245), .Z(n3344_adj_2043)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2202_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i31854_2_lut_4_lut (.A(n38293), .B(n4540[17]), .C(n38307), .D(n35898), 
         .Z(n36690)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i31854_2_lut_4_lut.init = 16'hffca;
    LUT4 i32078_4_lut (.A(n38397), .B(n38396), .C(n38400), .D(n36899), 
         .Z(n36914)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32078_4_lut.init = 16'h0100;
    LUT4 i32063_4_lut (.A(n38399), .B(n38376), .C(n38375), .D(n36886), 
         .Z(n36899)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32063_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_adj_337 (.A(n1709[27]), .B(n1709[28]), .Z(n34956)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_adj_337.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_338 (.A(n2342_adj_1771), .B(n2402_adj_2195[25]), 
         .C(n38267), .D(n2444_adj_1604), .Z(n36268)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_338.init = 16'hffca;
    LUT4 i32050_4_lut (.A(n38373), .B(n38395), .C(n38357), .D(n5_adj_2121), 
         .Z(n36886)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam i32050_4_lut.init = 16'h5554;
    CCU2C rem_10_add_2249_23 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[23]), 
          .D0(n3235_adj_539), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[24]), 
          .D1(n3234_adj_630), .CIN(n31118), .COUT(n31119), .S0(n3392_adj_2163[23]), 
          .S1(n3392_adj_2163[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_23.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_23.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_23.INJECT1_0 = "NO";
    defparam rem_10_add_2249_23.INJECT1_1 = "NO";
    CCU2C rem_10_add_2249_21 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[21]), 
          .D0(n3237_adj_542), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[22]), 
          .D1(n3236_adj_568), .CIN(n31117), .COUT(n31118), .S0(n3392_adj_2163[21]), 
          .S1(n3392_adj_2163[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_21.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_21.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_21.INJECT1_0 = "NO";
    defparam rem_10_add_2249_21.INJECT1_1 = "NO";
    LUT4 div_9_i2186_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[29]), 
         .D(n38190), .Z(n3328_adj_2044)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2186_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24360_2_lut_rep_262 (.A(n28297), .B(n13555), .Z(n38267)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24360_2_lut_rep_262.init = 16'heeee;
    LUT4 pwm_cnt_14__I_0_51_i5_2_lut (.A(pwm_cnt[2]), .B(duty3[2]), .Z(n5_adj_2121)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(104[20:37])
    defparam pwm_cnt_14__I_0_51_i5_2_lut.init = 16'h6666;
    LUT4 i32021_4_lut (.A(n38391), .B(n38390), .C(n38394), .D(n36842), 
         .Z(n36857)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32021_4_lut.init = 16'h0100;
    LUT4 div_9_i1587_3_lut_rep_261_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[25]), 
         .D(n2342_adj_1771), .Z(n38266)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1587_3_lut_rep_261_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut (.A(n3152), .B(n38202), .C(n3150), .Z(n33434)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 div_9_i1585_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[27]), 
         .D(n2340_adj_1746), .Z(n2439_adj_1317)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1585_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i23_3_lut (.A(n75_adj_8), .B(n38[22]), .C(n3556), 
         .Z(n329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i23_3_lut.init = 16'hcaca;
    LUT4 div_9_i1581_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[31]), 
         .D(n2336_adj_1708), .Z(n2435)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1581_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32006_4_lut (.A(n38393), .B(n38372), .C(n38371), .D(n36829), 
         .Z(n36842)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i32006_4_lut.init = 16'h5455;
    LUT4 div_9_i1599_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[13]), 
         .D(n2354_adj_1910), .Z(n2453_adj_1327)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1599_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2249_19 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[19]), 
          .D0(n3239_adj_624), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[20]), 
          .D1(n3238_adj_639), .CIN(n31116), .COUT(n31117), .S0(n3392_adj_2163[19]), 
          .S1(n3392_adj_2163[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_19.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_19.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_19.INJECT1_0 = "NO";
    defparam rem_10_add_2249_19.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_339 (.A(n34880), .B(n34790), .C(n1750_adj_1443), 
         .D(n28098), .Z(n28566)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_339.init = 16'ha8a0;
    LUT4 div_9_i1594_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[18]), 
         .D(n2349_adj_1861), .Z(n2448_adj_1321)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1594_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_340 (.A(n1748_adj_1438), .B(n1747_adj_1430), .C(n1749_adj_1436), 
         .Z(n34880)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_340.init = 16'h8080;
    LUT4 div_9_i1584_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[28]), 
         .D(n2339_adj_1739), .Z(n2438_adj_1312)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1584_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i31993_4_lut (.A(n38369), .B(n38389), .C(n38356), .D(n5_adj_2122), 
         .Z(n36829)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam i31993_4_lut.init = 16'h5554;
    LUT4 div_9_i1596_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[16]), 
         .D(n2351_adj_1867), .Z(n2450_adj_1324)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1596_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_341 (.A(n27382), .B(n3), .C(n45), .Z(duty0_14__N_426[13])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_341.init = 16'h2020;
    LUT4 pwm_cnt_14__I_0_52_i5_2_lut (.A(pwm_cnt[2]), .B(duty2[2]), .Z(n5_adj_2122)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(103[20:37])
    defparam pwm_cnt_14__I_0_52_i5_2_lut.init = 16'h6666;
    LUT4 i24147_3_lut (.A(n333_adj_1452), .B(n1753_adj_724), .C(n1754_adj_1454), 
         .Z(n28098)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24147_3_lut.init = 16'hecec;
    CCU2C rem_10_add_2249_17 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[17]), 
          .D0(n3241), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[18]), 
          .D1(n3240_adj_561), .CIN(n31115), .COUT(n31116), .S0(n3392_adj_2163[17]), 
          .S1(n3392_adj_2163[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_17.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_17.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_17.INJECT1_0 = "NO";
    defparam rem_10_add_2249_17.INJECT1_1 = "NO";
    LUT4 i31964_4_lut (.A(n38385), .B(n38384), .C(n38388), .D(n36785), 
         .Z(n36800)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i31964_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_342 (.A(n1742_adj_1423), .B(n35728), .C(n1746_adj_1432), 
         .D(n1745_adj_1425), .Z(n13638)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_342.init = 16'hfffe;
    LUT4 i31949_4_lut (.A(n38387), .B(n38368), .C(n38367), .D(n36772), 
         .Z(n36785)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i31949_4_lut.init = 16'h5455;
    LUT4 i1_2_lut_4_lut_adj_343 (.A(n3044), .B(n3095[16]), .C(n38204), 
         .D(n3133_adj_2014), .Z(n36056)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_343.init = 16'hffca;
    LUT4 i31936_4_lut (.A(n38365), .B(n38383), .C(n38355), .D(n5_adj_2123), 
         .Z(n36772)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam i31936_4_lut.init = 16'h5554;
    LUT4 pwm_cnt_14__I_0_53_i5_2_lut (.A(pwm_cnt[2]), .B(duty1[2]), .Z(n5_adj_2123)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(102[20:37])
    defparam pwm_cnt_14__I_0_53_i5_2_lut.init = 16'h6666;
    LUT4 div_9_i1600_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[12]), 
         .D(n339_adj_1752), .Z(n2454_adj_1328)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1600_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1583_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[29]), 
         .D(n2338_adj_1741), .Z(n2437_adj_1310)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1583_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21_4_lut (.A(n72_adj_5), .B(n38[28]), .C(n3556), .D(n38[23]), 
         .Z(n1354)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i21_4_lut.init = 16'h3aca;
    LUT4 i31907_4_lut (.A(n38379), .B(n38378), .C(n38382), .D(n36728), 
         .Z(n36743)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i31907_4_lut.init = 16'h0100;
    LUT4 div_9_i1593_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[19]), 
         .D(n2348_adj_1863), .Z(n2447_adj_1320)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1593_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i31892_4_lut (.A(n38381), .B(n38364), .C(n38363), .D(n36715), 
         .Z(n36728)) /* synthesis lut_function=(!(A+!(B+(C+!(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i31892_4_lut.init = 16'h5455;
    LUT4 div_9_i1592_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[20]), 
         .D(n2347_adj_1830), .Z(n2446_adj_1313)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1592_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i31879_4_lut (.A(n38361), .B(n38377), .C(n38354), .D(n5_adj_2124), 
         .Z(n36715)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam i31879_4_lut.init = 16'h5554;
    LUT4 div_9_i2193_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[22]), 
         .D(n3236), .Z(n3335_adj_1716)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2193_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_195_4_lut (.A(n3052), .B(n3095[8]), .C(n38204), 
         .D(n3152), .Z(n38200)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_rep_195_4_lut.init = 16'hca00;
    LUT4 pwm_cnt_14__I_0_54_i5_2_lut (.A(pwm_cnt[2]), .B(duty0[2]), .Z(n5_adj_2124)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(101[20:37])
    defparam pwm_cnt_14__I_0_54_i5_2_lut.init = 16'h6666;
    LUT4 select_842_Select_0_i4_3_lut_4_lut (.A(n38163), .B(n1), .C(n197[0]), 
         .D(n2983), .Z(duty0_14__N_410[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam select_842_Select_0_i4_3_lut_4_lut.init = 16'hff10;
    CCU2C rem_10_add_2249_15 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[15]), 
          .D0(n3243_adj_580), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[16]), 
          .D1(n3242_adj_588), .CIN(n31114), .COUT(n31115), .S0(n3392_adj_2163[15]), 
          .S1(n3392_adj_2163[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_15.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_15.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_15.INJECT1_0 = "NO";
    defparam rem_10_add_2249_15.INJECT1_1 = "NO";
    CCU2C rem_10_add_2249_13 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[13]), 
          .D0(n3245_adj_642), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[14]), 
          .D1(n3244_adj_551), .CIN(n31113), .COUT(n31114), .S0(n3392_adj_2163[13]), 
          .S1(n3392_adj_2163[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_13.INJECT1_0 = "NO";
    defparam rem_10_add_2249_13.INJECT1_1 = "NO";
    LUT4 div_9_i1597_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[15]), 
         .D(n2352_adj_1880), .Z(n2451_adj_1323)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1597_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_344 (.A(n1351), .B(n28391), .C(n1350), .D(n1448), 
         .Z(n28558)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_344.init = 16'h8000;
    LUT4 i24438_4_lut (.A(n28110), .B(n1352), .C(n1353), .D(n1354), 
         .Z(n28391)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24438_4_lut.init = 16'heccc;
    LUT4 i24159_3_lut (.A(n331), .B(n329), .C(n330), .Z(n28110)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24159_3_lut.init = 16'hecec;
    LUT4 div_9_i1591_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[21]), 
         .D(n38270), .Z(n2445_adj_1311)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1591_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i21_3_lut (.A(n81_adj_11), .B(n38[20]), .C(n3556), 
         .Z(n331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i21_3_lut.init = 16'hcaca;
    LUT4 div_13_mux_3_i22_3_lut (.A(n78_adj_7), .B(n38[21]), .C(n3556), 
         .Z(n330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i22_3_lut.init = 16'hcaca;
    LUT4 i26251_4_lut (.A(n66_adj_2), .B(n30240), .C(n38[25]), .D(n3556), 
         .Z(n6_adj_1495)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i26251_4_lut.init = 16'hfcee;
    LUT4 i26241_4_lut (.A(n69_adj_6), .B(n328), .C(n38[24]), .D(n3556), 
         .Z(n30240)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i26241_4_lut.init = 16'hc088;
    LUT4 div_9_i1586_3_lut_rep_260_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[26]), 
         .D(n2341_adj_1744), .Z(n38265)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1586_3_lut_rep_260_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i24_3_lut (.A(n72_adj_5), .B(n38[23]), .C(n3556), 
         .Z(n328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i24_3_lut.init = 16'hcaca;
    CCU2C rem_10_add_2249_11 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[11]), 
          .D0(n3247_adj_599), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[12]), 
          .D1(n3246), .CIN(n31112), .COUT(n31113), .S0(n3392_adj_2163[11]), 
          .S1(n3392_adj_2163[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_11.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_11.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_11.INJECT1_0 = "NO";
    defparam rem_10_add_2249_11.INJECT1_1 = "NO";
    LUT4 div_9_i1595_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[17]), 
         .D(n2350_adj_1869), .Z(n2449_adj_1322)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1595_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1589_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[23]), 
         .D(n2344_adj_1814), .Z(n2443_adj_1319)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1589_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1582_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[30]), 
         .D(n2337_adj_1706), .Z(n2436_adj_1318)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1582_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1590_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[22]), 
         .D(n2345_adj_1812), .Z(n2444_adj_1604)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1590_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1598_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[14]), 
         .D(n2353_adj_1878), .Z(n2452_adj_1325)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1598_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1588_3_lut_4_lut (.A(n28297), .B(n13555), .C(n2402_adj_2195[24]), 
         .D(n2343), .Z(n2442_adj_1601)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1588_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_345 (.A(n2238_adj_1833), .B(n2303_adj_2197[30]), 
         .C(n38269), .D(n2341_adj_1912), .Z(n35526)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_345.init = 16'hffca;
    LUT4 i24280_2_lut_rep_264 (.A(n28208), .B(n13616), .Z(n38269)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24280_2_lut_rep_264.init = 16'heeee;
    LUT4 rem_10_i1515_3_lut_rep_263_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[30]), 
         .D(n2238_adj_1833), .Z(n38268)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1515_3_lut_rep_263_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1523_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[22]), 
         .D(n2246_adj_1849), .Z(n2345_adj_1932)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1523_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_346 (.A(n2935_adj_2114), .B(n2996_adj_2201[26]), 
         .C(n38209), .D(n3040_adj_1116), .Z(n34988)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_346.init = 16'hffca;
    LUT4 i1_4_lut_adj_347 (.A(n31539), .B(n34948), .C(n34944), .D(n34942), 
         .Z(n27382)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_347.init = 16'hfffe;
    LUT4 i24628_2_lut_rep_199 (.A(n28578), .B(n13548), .Z(n38204)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24628_2_lut_rep_199.init = 16'heeee;
    LUT4 rem_10_i1529_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[16]), 
         .D(n2252_adj_1873), .Z(n2351_adj_1946)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1529_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1532_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[13]), 
         .D(n587), .Z(n2354_adj_1954)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1532_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2073_3_lut_rep_197_4_lut (.A(n28578), .B(n13548), .C(n3095[8]), 
         .D(n3052), .Z(n38202)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2073_3_lut_rep_197_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2050_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[31]), 
         .D(n3029), .Z(n3128_adj_1528)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2050_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2249_9 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[9]), 
          .D0(n3249_adj_622), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[10]), 
          .D1(n3248_adj_618), .CIN(n31111), .COUT(n31112), .S0(n3392_adj_2163[9]), 
          .S1(n3392_adj_2163[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_9.INIT0 = 16'hf1e0;
    defparam rem_10_add_2249_9.INIT1 = 16'hf1e0;
    defparam rem_10_add_2249_9.INJECT1_0 = "NO";
    defparam rem_10_add_2249_9.INJECT1_1 = "NO";
    CCU2C rem_10_add_2249_7 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[7]), 
          .D0(n3251), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[8]), 
          .D1(n3250), .CIN(n31110), .COUT(n31111), .S0(n3392_adj_2163[7]), 
          .S1(n3392_adj_2163[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_7.INIT0 = 16'h0e1f;
    defparam rem_10_add_2249_7.INIT1 = 16'hf1e0;
    defparam rem_10_add_2249_7.INJECT1_0 = "NO";
    defparam rem_10_add_2249_7.INJECT1_1 = "NO";
    LUT4 rem_10_i1526_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[19]), 
         .D(n2249_adj_1852), .Z(n2348_adj_1943)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1526_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1514_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[31]), 
         .D(n2237_adj_1827), .Z(n2336_adj_1900)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1514_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1516_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[29]), 
         .D(n2239_adj_1832), .Z(n2338_adj_1905)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1516_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1522_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[23]), 
         .D(n2245_adj_1844), .Z(n2344_adj_1933)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1522_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1528_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[17]), 
         .D(n2251_adj_1856), .Z(n2350_adj_1947)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1528_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2195_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[20]), 
         .D(n3238), .Z(n3337_adj_1526)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2195_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1517_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[28]), 
         .D(n2240_adj_1837), .Z(n2339_adj_1904)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1517_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2066_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[15]), 
         .D(n3045), .Z(n3144)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2066_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2249_5 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[5]), 
          .D0(n3253_adj_1776), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[6]), 
          .D1(n38198), .CIN(n31109), .COUT(n31110), .S0(n3392_adj_2163[5]), 
          .S1(n3392_adj_2163[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_5.INIT0 = 16'hf1e0;
    defparam rem_10_add_2249_5.INIT1 = 16'hf1e0;
    defparam rem_10_add_2249_5.INJECT1_0 = "NO";
    defparam rem_10_add_2249_5.INJECT1_1 = "NO";
    LUT4 div_13_mux_3_i16_3_lut (.A(n96), .B(n38[15]), .C(n3556), .Z(n336_adj_1064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i16_3_lut.init = 16'hcaca;
    CCU2C rem_10_add_2249_3 (.A0(n13620), .B0(n28434), .C0(n3293_adj_2161[3]), 
          .D0(n597), .A1(n13620), .B1(n28434), .C1(n3293_adj_2161[4]), 
          .D1(n3254_adj_597), .CIN(n31108), .COUT(n31109), .S0(n3392_adj_2163[3]), 
          .S1(n3392_adj_2163[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_3.INIT0 = 16'hf1e0;
    defparam rem_10_add_2249_3.INIT1 = 16'h0e1f;
    defparam rem_10_add_2249_3.INJECT1_0 = "NO";
    defparam rem_10_add_2249_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1518_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[27]), 
         .D(n2241_adj_1836), .Z(n2340_adj_1913)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1518_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2249_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(distance[0]), .D1(n2[2]), 
          .COUT(n31108), .S1(n3392_adj_2163[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2249_1.INIT0 = 16'h0000;
    defparam rem_10_add_2249_1.INIT1 = 16'habef;
    defparam rem_10_add_2249_1.INJECT1_0 = "NO";
    defparam rem_10_add_2249_1.INJECT1_1 = "NO";
    LUT4 div_9_i2056_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[25]), 
         .D(n3035), .Z(n3134)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2056_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2059_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[22]), 
         .D(n3038), .Z(n3137)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2059_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2361_12 (.A0(n3545), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n31107), .S0(n3568[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2361_12.INIT0 = 16'h5550;
    defparam rem_10_add_2361_12.INIT1 = 16'h0000;
    defparam rem_10_add_2361_12.INJECT1_0 = "NO";
    defparam rem_10_add_2361_12.INJECT1_1 = "NO";
    CCU2C rem_10_add_2361_10 (.A0(n3547), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n3546), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31106), .COUT(n31107), .S0(n3568[8]), .S1(n3568[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2361_10.INIT0 = 16'h5550;
    defparam rem_10_add_2361_10.INIT1 = 16'h5550;
    defparam rem_10_add_2361_10.INJECT1_0 = "NO";
    defparam rem_10_add_2361_10.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_348 (.A(n1709[29]), .B(n1709[30]), .Z(n34958)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_adj_348.init = 16'heeee;
    LUT4 div_9_i2201_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[14]), 
         .D(n3244), .Z(n3343_adj_1525)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2201_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2076_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[5]), 
         .D(n346), .Z(n3154)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2076_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1520_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[25]), 
         .D(n2243_adj_1840), .Z(n2342_adj_1929)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1520_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i3_3_lut (.A(n135), .B(n38[2]), .C(n3556), .Z(n349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i3_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1527_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[18]), 
         .D(n2250_adj_1857), .Z(n2349_adj_1942)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1527_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i4_3_lut (.A(n132), .B(n38[3]), .C(n3556), .Z(n348_adj_1735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i4_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1525_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[20]), 
         .D(n2248_adj_1853), .Z(n2347_adj_1936)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1525_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1524_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[21]), 
         .D(n2247_adj_1848), .Z(n2346_adj_1937)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1524_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i5_3_lut (.A(n129), .B(n38[4]), .C(n3556), .Z(n347_adj_667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i5_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1519_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[26]), 
         .D(n2242_adj_1841), .Z(n2341_adj_1912)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1519_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1521_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[24]), 
         .D(n2244_adj_1845), .Z(n2343_adj_1928)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1521_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1531_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[14]), 
         .D(n2254_adj_1889), .Z(n2353_adj_1950)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1531_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i7_3_lut (.A(n123), .B(n38[6]), .C(n3556), .Z(n345_adj_2111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i7_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1530_3_lut_4_lut (.A(n28208), .B(n13616), .C(n2303_adj_2197[15]), 
         .D(n2253_adj_1872), .Z(n2352_adj_1951)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i1530_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2361_8 (.A0(n3549), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n3548), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31105), 
          .COUT(n31106), .S0(n3568[6]), .S1(n3568[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2361_8.INIT0 = 16'h5550;
    defparam rem_10_add_2361_8.INIT1 = 16'h5550;
    defparam rem_10_add_2361_8.INJECT1_0 = "NO";
    defparam rem_10_add_2361_8.INJECT1_1 = "NO";
    CCU2C rem_10_add_2361_6 (.A0(n3551), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n3550), .B1(GND_net), .C1(GND_net), .D1(VCC_net), .CIN(n31104), 
          .COUT(n31105), .S0(n3568[4]), .S1(n3568[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2361_6.INIT0 = 16'h5550;
    defparam rem_10_add_2361_6.INIT1 = 16'h5550;
    defparam rem_10_add_2361_6.INJECT1_0 = "NO";
    defparam rem_10_add_2361_6.INJECT1_1 = "NO";
    LUT4 div_13_i1452_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[26]), 
         .D(n2143_adj_984), .Z(n2242)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1452_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i6_3_lut (.A(n126), .B(n38[5]), .C(n3556), .Z(n346_adj_1140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i6_3_lut.init = 16'hcaca;
    LUT4 div_13_i1458_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[20]), 
         .D(n2149_adj_994), .Z(n2248)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1458_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2051_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[30]), 
         .D(n38212), .Z(n3129)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2051_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1451_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[27]), 
         .D(n2142_adj_990), .Z(n2241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1451_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2361_4 (.A0(n3454), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n3453), .B1(n3458), .C1(GND_net), .D1(VCC_net), .CIN(n31103), 
          .COUT(n31104), .S0(n3568[2]), .S1(n3568[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2361_4.INIT0 = 16'h5550;
    defparam rem_10_add_2361_4.INIT1 = 16'h9999;
    defparam rem_10_add_2361_4.INJECT1_0 = "NO";
    defparam rem_10_add_2361_4.INJECT1_1 = "NO";
    LUT4 div_13_i2405_3_lut_4_lut (.A(n28412), .B(n13634), .C(n3556), 
         .D(n4990[13]), .Z(n197[13])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i2405_3_lut_4_lut.init = 16'hfe0e;
    LUT4 div_9_i2065_3_lut_rep_196_4_lut (.A(n28578), .B(n13548), .C(n3095[16]), 
         .D(n3044), .Z(n38201)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2065_3_lut_rep_196_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1462_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[16]), 
         .D(n2153_adj_1002), .Z(n2252)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1462_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1449_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[29]), 
         .D(n2140_adj_991), .Z(n2239)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1449_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_add_2361_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n33580), .B1(n33697), .C1(GND_net), .D1(VCC_net), 
          .COUT(n31103), .S1(n3568[1]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_2361_2.INIT0 = 16'h000f;
    defparam rem_10_add_2361_2.INIT1 = 16'h1111;
    defparam rem_10_add_2361_2.INJECT1_0 = "NO";
    defparam rem_10_add_2361_2.INJECT1_1 = "NO";
    LUT4 div_9_i2061_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[20]), 
         .D(n3040), .Z(n3139)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2061_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1460_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[18]), 
         .D(n2151_adj_995), .Z(n2250)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1460_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i11_3_lut (.A(n111), .B(n38[10]), .C(n3556), .Z(n341_adj_605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i11_3_lut.init = 16'hcaca;
    PFUMX i32320 (.BLUT(n37671), .ALUT(n37670), .C0(n38177), .Z(n37672));
    LUT4 div_13_i1461_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[17]), 
         .D(n2152), .Z(n2251)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1461_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1457_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[21]), 
         .D(n2148_adj_992), .Z(n2247)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1457_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1456_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[22]), 
         .D(n2147_adj_993), .Z(n2246)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1456_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1463_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[15]), 
         .D(n2154_adj_1003), .Z(n2253)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1463_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1454_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[24]), 
         .D(n2145), .Z(n2244)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1454_3_lut_4_lut.init = 16'hf1e0;
    CCU2C pwm_cnt_1138_add_4_15 (.A0(pwm_cnt[13]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[14]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31101), .S0(n50[13]), .S1(n50[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_15.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_15.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_15.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_15.INJECT1_1 = "NO";
    CCU2C pwm_cnt_1138_add_4_13 (.A0(pwm_cnt[11]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[12]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31100), .COUT(n31101), .S0(n50[11]), .S1(n50[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_13.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_13.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_13.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_13.INJECT1_1 = "NO";
    LUT4 div_9_i2057_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[24]), 
         .D(n3036), .Z(n3135)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2057_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1450_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[28]), 
         .D(n2141_adj_983), .Z(n2240)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1450_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1447_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[31]), 
         .D(n2138), .Z(n2237)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1447_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1448_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[30]), 
         .D(n2139), .Z(n2238)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1448_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1459_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[19]), 
         .D(n2150_adj_996), .Z(n2249)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1459_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1464_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[14]), 
         .D(n337_adj_1001), .Z(n2254)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1464_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1453_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[25]), 
         .D(n2144_adj_986), .Z(n2243)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1453_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i9_3_lut (.A(n117), .B(n38[8]), .C(n3556), .Z(n343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i9_3_lut.init = 16'hcaca;
    LUT4 div_13_i1455_3_lut_4_lut (.A(n28412), .B(n13634), .C(n2204_adj_2174[23]), 
         .D(n2146_adj_985), .Z(n2245)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1455_3_lut_4_lut.init = 16'hf1e0;
    CCU2C pwm_cnt_1138_add_4_11 (.A0(pwm_cnt[9]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[10]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31099), .COUT(n31100), .S0(n50[9]), .S1(n50[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_11.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_11.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_11.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_349 (.A(n2247_adj_2017), .B(n2303[21]), .C(n38271), 
         .D(n2343), .Z(n36234)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_349.init = 16'hffca;
    LUT4 i24322_2_lut_rep_266 (.A(n28269), .B(n13557), .Z(n38271)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24322_2_lut_rep_266.init = 16'heeee;
    LUT4 div_9_i1524_3_lut_rep_265_4_lut (.A(n28269), .B(n13557), .C(n2303[21]), 
         .D(n2247_adj_2017), .Z(n38270)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1524_3_lut_rep_265_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1529_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[16]), 
         .D(n2252_adj_2091), .Z(n2351_adj_1867)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1529_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1528_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[17]), 
         .D(n2251_adj_2089), .Z(n2350_adj_1869)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1528_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1523_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[22]), 
         .D(n2246_adj_2018), .Z(n2345_adj_1812)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1523_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i10_3_lut (.A(n114), .B(n38[9]), .C(n3556), .Z(n342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i10_3_lut.init = 16'hcaca;
    LUT4 div_9_i2190_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[25]), 
         .D(n3233_adj_522), .Z(n3332_adj_1527)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1522_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[23]), 
         .D(n2245_adj_2015), .Z(n2344_adj_1814)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1522_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2053_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[28]), 
         .D(n3032), .Z(n3131_adj_1727)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2053_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1518_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[27]), 
         .D(n2241_adj_1921), .Z(n2340_adj_1746)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1518_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1526_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[19]), 
         .D(n2249_adj_2087), .Z(n2348_adj_1863)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1526_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1519_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[26]), 
         .D(n2242_adj_1925), .Z(n2341_adj_1744)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1519_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1530_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[15]), 
         .D(n2253_adj_2092), .Z(n2352_adj_1880)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1530_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1527_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[18]), 
         .D(n2250_adj_2090), .Z(n2349_adj_1861)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1527_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_350 (.A(n36316), .B(n36318), .C(n36310), .D(n36314), 
         .Z(n13590)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_4_lut_adj_350.init = 16'hfffe;
    LUT4 i1_3_lut_adj_351 (.A(n2142), .B(n2146), .C(n2144), .Z(n36318)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_3_lut_adj_351.init = 16'hfefe;
    LUT4 i1_4_lut_adj_352 (.A(n35930), .B(n35784), .C(n2150), .D(n27984), 
         .Z(n28440)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_352.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_353 (.A(n2147), .B(n2148), .C(n2149), .Z(n35930)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_353.init = 16'h8080;
    CCU2C pwm_cnt_1138_add_4_9 (.A0(pwm_cnt[7]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[8]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31098), .COUT(n31099), .S0(n50[7]), .S1(n50[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_9.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_9.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_9.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_9.INJECT1_1 = "NO";
    CCU2C pwm_cnt_1138_add_4_7 (.A0(pwm_cnt[5]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[6]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31097), .COUT(n31098), .S0(n50[5]), .S1(n50[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_7.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_7.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_7.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_7.INJECT1_1 = "NO";
    LUT4 i24034_3_lut (.A(n337), .B(n2153), .C(n2154), .Z(n27984)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24034_3_lut.init = 16'hecec;
    LUT4 div_9_i1532_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[13]), 
         .D(n338), .Z(n2354_adj_1910)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1532_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1516_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[29]), 
         .D(n2239_adj_1917), .Z(n2338_adj_1741)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1516_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1517_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[28]), 
         .D(n2240_adj_1922), .Z(n2339_adj_1739)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1517_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1525_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[20]), 
         .D(n2248_adj_2086), .Z(n2347_adj_1830)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1525_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2406_3_lut_rep_161_4_lut (.A(n28269), .B(n13557), .C(n38307), 
         .D(n4540[12]), .Z(n38166)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_9_i2406_3_lut_rep_161_4_lut.init = 16'hfe0e;
    CCU2C pwm_cnt_1138_add_4_5 (.A0(pwm_cnt[3]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[4]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31096), .COUT(n31097), .S0(n50[3]), .S1(n50[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_5.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_5.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_5.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_5.INJECT1_1 = "NO";
    CCU2C pwm_cnt_1138_add_4_3 (.A0(pwm_cnt[1]), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(pwm_cnt[2]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .CIN(n31095), .COUT(n31096), .S0(n50[1]), .S1(n50[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_3.INIT0 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_3.INIT1 = 16'haaa0;
    defparam pwm_cnt_1138_add_4_3.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_3.INJECT1_1 = "NO";
    LUT4 div_9_i1514_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[31]), 
         .D(n2237_adj_1916), .Z(n2336_adj_1708)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1514_3_lut_4_lut.init = 16'hf1e0;
    CCU2C pwm_cnt_1138_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_cnt[0]), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n31095), .S1(n50[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(96[23:37])
    defparam pwm_cnt_1138_add_4_1.INIT0 = 16'h0000;
    defparam pwm_cnt_1138_add_4_1.INIT1 = 16'h555f;
    defparam pwm_cnt_1138_add_4_1.INJECT1_0 = "NO";
    defparam pwm_cnt_1138_add_4_1.INJECT1_1 = "NO";
    CCU2C div_9_unary_minus_2_add_3_19 (.A0(n5), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n31094), .S0(n35[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_19.INIT0 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_19.INIT1 = 16'h0000;
    defparam div_9_unary_minus_2_add_3_19.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_19.INJECT1_1 = "NO";
    LUT4 i28743_2_lut (.A(n1610[29]), .B(n28558), .Z(n1645)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i28743_2_lut.init = 16'h8888;
    LUT4 div_9_i1520_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[25]), 
         .D(n2243_adj_1924), .Z(n2342_adj_1771)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1520_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_unary_minus_2_add_3_17 (.A0(n39), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n5), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31093), .COUT(n31094), .S0(n35[17]), .S1(n35[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_17.INIT0 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_17.INIT1 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_17.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_17.INJECT1_1 = "NO";
    LUT4 div_9_i1515_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[30]), 
         .D(n2238_adj_1918), .Z(n2337_adj_1706)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1515_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1521_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[24]), 
         .D(n2244_adj_2016), .Z(n2343)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1521_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_unary_minus_2_add_3_15 (.A0(n45), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n42), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31092), .COUT(n31093), .S0(n35[15]), .S1(n35[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_15.INIT0 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_15.INIT1 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_15.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_15.INJECT1_1 = "NO";
    LUT4 div_9_i2068_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[13]), 
         .D(n3047), .Z(n3146)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2068_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1531_3_lut_4_lut (.A(n28269), .B(n13557), .C(n2303[14]), 
         .D(n2254_adj_2093), .Z(n2353_adj_1878)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i1531_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2074_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[7]), 
         .D(n3053), .Z(n3152)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2074_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i28736_2_lut (.A(n1610[31]), .B(n28558), .Z(n1643)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i28736_2_lut.init = 16'h8888;
    LUT4 div_13_i1385_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[26]), 
         .D(n2044_adj_1050), .Z(n2143_adj_984)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1385_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2203_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[12]), 
         .D(n3246_adj_548), .Z(n3345_adj_1715)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2203_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2404_3_lut_4_lut (.A(n28401), .B(n13635), .C(n3556), 
         .D(n4990[14]), .Z(n197[14])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i2404_3_lut_4_lut.init = 16'hfe0e;
    CCU2C div_9_unary_minus_2_add_3_13 (.A0(n51), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n48), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31091), .COUT(n31092), .S0(n35[13]), .S1(n35[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_13.INIT0 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_13.INIT1 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_13.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_13.INJECT1_1 = "NO";
    CCU2C div_9_unary_minus_2_add_3_11 (.A0(n38317), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n54), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31090), .COUT(n31091), .S0(n35[11]), .S1(n35[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_11.INIT0 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_11.INIT1 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_11.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_11.INJECT1_1 = "NO";
    LUT4 div_13_i1383_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[28]), 
         .D(n2042_adj_1053), .Z(n2141_adj_983)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1383_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1391_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[20]), 
         .D(n2050_adj_1062), .Z(n2149_adj_994)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1391_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1381_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[30]), 
         .D(n2040_adj_1051), .Z(n2139)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1381_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_unary_minus_2_add_3_9 (.A0(n38322), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n38316), .B1(n27382), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31089), .COUT(n31090), .S0(n35[9]), .S1(n35[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_9.INIT0 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_9.INIT1 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_9.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_9.INJECT1_1 = "NO";
    LUT4 div_13_i1384_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[27]), 
         .D(n2043_adj_1049), .Z(n2142_adj_990)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1384_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_unary_minus_2_add_3_7 (.A0(n38332), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n66_adj_9), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31088), .COUT(n31089), .S0(n35[7]), .S1(n35[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_7.INIT0 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_7.INIT1 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_7.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_7.INJECT1_1 = "NO";
    LUT4 div_9_i2062_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[19]), 
         .D(n3041), .Z(n3140)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2062_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_9_unary_minus_2_add_3_5 (.A0(n75_adj_1), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n38333), .B1(n27382), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31087), .COUT(n31088), .S0(n35[5]), .S1(n35[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_5.INIT0 = 16'hdddd;
    defparam div_9_unary_minus_2_add_3_5.INIT1 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_5.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_5.INJECT1_1 = "NO";
    CCU2C div_9_unary_minus_2_add_3_3 (.A0(n38335), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n38334), .B1(n27382), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31086), .COUT(n31087), .S0(n35[3]), .S1(n35[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_3.INIT0 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_3.INIT1 = 16'h7777;
    defparam div_9_unary_minus_2_add_3_3.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_3.INJECT1_1 = "NO";
    CCU2C div_9_unary_minus_2_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[0]), .B1(n12154), .C1(GND_net), 
          .D1(VCC_net), .COUT(n31086), .S1(n35[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_unary_minus_2_add_3_1.INIT0 = 16'h0000;
    defparam div_9_unary_minus_2_add_3_1.INIT1 = 16'h222d;
    defparam div_9_unary_minus_2_add_3_1.INJECT1_0 = "NO";
    defparam div_9_unary_minus_2_add_3_1.INJECT1_1 = "NO";
    CCU2C rem_10_unary_minus_2_add_3_19 (.A0(n5), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n31085), .S0(n2[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_19.INIT0 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_19.INIT1 = 16'h0000;
    defparam rem_10_unary_minus_2_add_3_19.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_19.INJECT1_1 = "NO";
    CCU2C rem_10_unary_minus_2_add_3_17 (.A0(n39), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n5), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31084), .COUT(n31085), .S0(n2[17]), .S1(n2[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_17.INIT0 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_17.INIT1 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_17.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_17.INJECT1_1 = "NO";
    CCU2C rem_10_unary_minus_2_add_3_15 (.A0(n45), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n42), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31083), .COUT(n31084), .S0(n2[15]), .S1(n2[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_15.INIT0 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_15.INIT1 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_15.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_15.INJECT1_1 = "NO";
    LUT4 div_13_i1395_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[16]), 
         .D(n2054_adj_1066), .Z(n2153_adj_1002)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1395_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1386_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[25]), 
         .D(n2045_adj_1048), .Z(n2144_adj_986)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1386_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1387_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[24]), 
         .D(n2046_adj_1052), .Z(n2145)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1387_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_unary_minus_2_add_3_13 (.A0(n51), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n48), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31082), .COUT(n31083), .S0(n2[13]), .S1(n2[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_13.INIT0 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_13.INIT1 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_13.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_13.INJECT1_1 = "NO";
    LUT4 div_13_mux_3_i19_3_lut (.A(n87), .B(n38[18]), .C(n3556), .Z(n333_adj_1452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i19_3_lut.init = 16'hcaca;
    LUT4 div_13_i1389_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[22]), 
         .D(n2048_adj_1058), .Z(n2147_adj_993)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1389_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1396_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[15]), 
         .D(n336_adj_1064), .Z(n2154_adj_1003)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1396_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_unary_minus_2_add_3_11 (.A0(n38317), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n54), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31081), .COUT(n31082), .S0(n2[11]), .S1(n2[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_11.INIT0 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_11.INIT1 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_11.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_354 (.A(n34774), .B(n34772), .C(distance[0]), .D(distance[1]), 
         .Z(n31539)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_354.init = 16'ha888;
    CCU2C rem_10_unary_minus_2_add_3_9 (.A0(n38322), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n38316), .B1(n27382), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31080), .COUT(n31081), .S0(n2[9]), .S1(n2[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_9.INIT0 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_9.INIT1 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_9.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_9.INJECT1_1 = "NO";
    LUT4 div_9_i2070_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[11]), 
         .D(n3049), .Z(n3148)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2070_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2052_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[29]), 
         .D(n38211), .Z(n3130)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2052_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_unary_minus_2_add_3_7 (.A0(n38332), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n66_adj_9), .B1(n12154), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31079), .COUT(n31080), .S0(n2[7]), .S1(n2[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_7.INIT0 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_7.INIT1 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_7.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_7.INJECT1_1 = "NO";
    LUT4 div_13_i1394_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[17]), 
         .D(n2053_adj_1065), .Z(n2152)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1394_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1382_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[29]), 
         .D(n2041_adj_1109), .Z(n2140_adj_991)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1382_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1380_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[31]), 
         .D(n38273), .Z(n2138)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1380_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1393_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[18]), 
         .D(n2052_adj_1063), .Z(n2151_adj_995)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1393_3_lut_4_lut.init = 16'hf1e0;
    CCU2C rem_10_unary_minus_2_add_3_5 (.A0(n75_adj_1), .B0(n12154), .C0(GND_net), 
          .D0(VCC_net), .A1(n38333), .B1(n27382), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31078), .COUT(n31079), .S0(n2[5]), .S1(n2[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_5.INIT0 = 16'hdddd;
    defparam rem_10_unary_minus_2_add_3_5.INIT1 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_5.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_5.INJECT1_1 = "NO";
    CCU2C rem_10_unary_minus_2_add_3_3 (.A0(n38335), .B0(n27382), .C0(GND_net), 
          .D0(VCC_net), .A1(n38334), .B1(n27382), .C1(GND_net), .D1(VCC_net), 
          .CIN(n31077), .COUT(n31078), .S0(n2[3]), .S1(n2[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_3.INIT0 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_3.INIT1 = 16'h7777;
    defparam rem_10_unary_minus_2_add_3_3.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_3.INJECT1_1 = "NO";
    CCU2C rem_10_unary_minus_2_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(distance[0]), .B1(n12154), .C1(GND_net), 
          .D1(VCC_net), .COUT(n31077), .S1(n2[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_unary_minus_2_add_3_1.INIT0 = 16'h0000;
    defparam rem_10_unary_minus_2_add_3_1.INIT1 = 16'h222d;
    defparam rem_10_unary_minus_2_add_3_1.INJECT1_0 = "NO";
    defparam rem_10_unary_minus_2_add_3_1.INJECT1_1 = "NO";
    LUT4 div_13_i1390_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[21]), 
         .D(n2049_adj_1060), .Z(n2148_adj_992)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1390_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2069_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[12]), 
         .D(n3048), .Z(n3147)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2069_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1388_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[23]), 
         .D(n2047_adj_1059), .Z(n2146_adj_985)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1388_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_1455_15 (.A0(n28412), .B0(n13634), .C0(GND_net), .D0(VCC_net), 
          .A1(n28401), .B1(n13635), .C1(GND_net), .D1(VCC_net), .CIN(n31075), 
          .S0(n4990[13]), .S1(n4990[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_15.INIT0 = 16'h1111;
    defparam add_1455_15.INIT1 = 16'h1111;
    defparam add_1455_15.INJECT1_0 = "NO";
    defparam add_1455_15.INJECT1_1 = "NO";
    CCU2C add_1455_13 (.A0(n28442), .B0(n13630), .C0(GND_net), .D0(VCC_net), 
          .A1(n28430), .B1(n13633), .C1(GND_net), .D1(VCC_net), .CIN(n31074), 
          .COUT(n31075), .S0(n4990[11]), .S1(n4990[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_13.INIT0 = 16'h1111;
    defparam add_1455_13.INIT1 = 16'h1111;
    defparam add_1455_13.INJECT1_0 = "NO";
    defparam add_1455_13.INJECT1_1 = "NO";
    CCU2C add_1455_11 (.A0(n28456), .B0(n13625), .C0(GND_net), .D0(VCC_net), 
          .A1(n28446), .B1(n13627), .C1(GND_net), .D1(VCC_net), .CIN(n31073), 
          .COUT(n31074), .S0(n4990[9]), .S1(n4990[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_11.INIT0 = 16'h1111;
    defparam add_1455_11.INIT1 = 16'h1111;
    defparam add_1455_11.INJECT1_0 = "NO";
    defparam add_1455_11.INJECT1_1 = "NO";
    LUT4 div_13_i1392_3_lut_4_lut (.A(n28401), .B(n13635), .C(n2105_adj_2178[19]), 
         .D(n2051_adj_1061), .Z(n2150_adj_996)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1392_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1461_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[17]), 
         .D(n2152_adj_1820), .Z(n2251_adj_1856)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1461_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2192_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[23]), 
         .D(n3235), .Z(n3334_adj_1714)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1462_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[16]), 
         .D(n2153_adj_1819), .Z(n2252_adj_1873)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1462_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2207_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[8]), 
         .D(n3250_adj_554), .Z(n3349_adj_2034)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2207_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i17_3_lut (.A(n93), .B(n38[16]), .C(n3556), .Z(n335_adj_1150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i17_3_lut.init = 16'hcaca;
    LUT4 rem_10_i1451_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[27]), 
         .D(n2142_adj_1794), .Z(n2241_adj_1836)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1451_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_1455_9 (.A0(n28468), .B0(n13622), .C0(GND_net), .D0(VCC_net), 
          .A1(n28462), .B1(n13624), .C1(GND_net), .D1(VCC_net), .CIN(n31072), 
          .COUT(n31073), .S0(n4990[7]), .S1(n4990[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_9.INIT0 = 16'h1111;
    defparam add_1455_9.INIT1 = 16'h1111;
    defparam add_1455_9.INJECT1_0 = "NO";
    defparam add_1455_9.INJECT1_1 = "NO";
    CCU2C add_1455_7 (.A0(n28506), .B0(n13618), .C0(GND_net), .D0(VCC_net), 
          .A1(n28484), .B1(n13621), .C1(GND_net), .D1(VCC_net), .CIN(n31071), 
          .COUT(n31072), .S0(n4990[5]), .S1(n4990[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_7.INIT0 = 16'h1111;
    defparam add_1455_7.INIT1 = 16'h1111;
    defparam add_1455_7.INJECT1_0 = "NO";
    defparam add_1455_7.INJECT1_1 = "NO";
    CCU2C add_1455_5 (.A0(n28522), .B0(n13614), .C0(GND_net), .D0(VCC_net), 
          .A1(n28518), .B1(n13617), .C1(GND_net), .D1(VCC_net), .CIN(n31070), 
          .COUT(n31071), .S0(n4990[3]), .S1(n4990[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_5.INIT0 = 16'h1111;
    defparam add_1455_5.INIT1 = 16'h1111;
    defparam add_1455_5.INJECT1_0 = "NO";
    defparam add_1455_5.INJECT1_1 = "NO";
    CCU2C add_1455_3 (.A0(n28267), .B0(n13608), .C0(GND_net), .D0(VCC_net), 
          .A1(n28528), .B1(n13610), .C1(GND_net), .D1(VCC_net), .CIN(n31069), 
          .COUT(n31070), .S0(n4990[1]), .S1(n4990[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_3.INIT0 = 16'h1111;
    defparam add_1455_3.INIT1 = 16'h1111;
    defparam add_1455_3.INJECT1_0 = "NO";
    defparam add_1455_3.INJECT1_1 = "NO";
    CCU2C add_1455_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n28303), .B1(n13607), .C1(GND_net), .D1(VCC_net), .COUT(n31069), 
          .S1(n4990[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam add_1455_1.INIT0 = 16'h0000;
    defparam add_1455_1.INIT1 = 16'heee1;
    defparam add_1455_1.INJECT1_0 = "NO";
    defparam add_1455_1.INJECT1_1 = "NO";
    LUT4 rem_10_i1459_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[19]), 
         .D(n2150_adj_1816), .Z(n2249_adj_1852)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1459_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2055_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[26]), 
         .D(n3034), .Z(n3133_adj_2014)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2055_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_31 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[31]), 
          .D0(n3227_adj_726), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31068), .S0(n3392_adj_2177[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_31.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_31.INIT1 = 16'h0000;
    defparam div_13_add_2249_31.INJECT1_0 = "NO";
    defparam div_13_add_2249_31.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_29 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[29]), 
          .D0(n3229_adj_723), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[30]), 
          .D1(n3228_adj_682), .CIN(n31067), .COUT(n31068), .S0(n3392_adj_2177[29]), 
          .S1(n3392_adj_2177[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_29.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_29.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_29.INJECT1_0 = "NO";
    defparam div_13_add_2249_29.INJECT1_1 = "NO";
    LUT4 rem_10_i1456_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[22]), 
         .D(n2147_adj_1803), .Z(n2246_adj_1849)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1456_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1447_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[31]), 
         .D(n2138_adj_1786), .Z(n2237_adj_1827)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1447_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_27 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[27]), 
          .D0(n3231_adj_612), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[28]), 
          .D1(n38182), .CIN(n31066), .COUT(n31067), .S0(n3392_adj_2177[27]), 
          .S1(n3392_adj_2177[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_27.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_27.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_27.INJECT1_0 = "NO";
    defparam div_13_add_2249_27.INJECT1_1 = "NO";
    LUT4 rem_10_i1460_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[18]), 
         .D(n2151_adj_1815), .Z(n2250_adj_1857)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1460_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2075_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[6]), 
         .D(n3054), .Z(n3153)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2075_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_25 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[25]), 
          .D0(n3233_adj_795), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[26]), 
          .D1(n3232_adj_766), .CIN(n31065), .COUT(n31066), .S0(n3392_adj_2177[25]), 
          .S1(n3392_adj_2177[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_25.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_25.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_25.INJECT1_0 = "NO";
    defparam div_13_add_2249_25.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_23 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[23]), 
          .D0(n3235_adj_792), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[24]), 
          .D1(n3234_adj_688), .CIN(n31064), .COUT(n31065), .S0(n3392_adj_2177[23]), 
          .S1(n3392_adj_2177[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_23.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_23.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_23.INJECT1_0 = "NO";
    defparam div_13_add_2249_23.INJECT1_1 = "NO";
    LUT4 div_9_i2205_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[10]), 
         .D(n3248), .Z(n3347_adj_1112)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2205_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_355 (.A(n38293), .B(n4540[17]), .C(n38307), 
         .D(n38166), .Z(n35902)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_355.init = 16'hffca;
    CCU2C div_13_add_2249_21 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[21]), 
          .D0(n3237_adj_662), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[22]), 
          .D1(n3236_adj_675), .CIN(n31063), .COUT(n31064), .S0(n3392_adj_2177[21]), 
          .S1(n3392_adj_2177[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_21.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_21.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_21.INJECT1_0 = "NO";
    defparam div_13_add_2249_21.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_19 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[19]), 
          .D0(n3239_adj_773), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[20]), 
          .D1(n3238_adj_754), .CIN(n31062), .COUT(n31063), .S0(n3392_adj_2177[19]), 
          .S1(n3392_adj_2177[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_19.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_19.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_19.INJECT1_0 = "NO";
    defparam div_13_add_2249_19.INJECT1_1 = "NO";
    LUT4 rem_10_i1450_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[28]), 
         .D(n2141_adj_1789), .Z(n2240_adj_1837)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1450_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2199_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[16]), 
         .D(n3242), .Z(n3341_adj_1114)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2199_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1453_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[25]), 
         .D(n2144_adj_1798), .Z(n2243_adj_1840)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1453_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2200_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[15]), 
         .D(n3243), .Z(n3342_adj_1713)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2200_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_17 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[17]), 
          .D0(n3241_adj_685), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[18]), 
          .D1(n3240_adj_564), .CIN(n31061), .COUT(n31062), .S0(n3392_adj_2177[17]), 
          .S1(n3392_adj_2177[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_17.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_17.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_17.INJECT1_0 = "NO";
    defparam div_13_add_2249_17.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_15 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[15]), 
          .D0(n3243_adj_692), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[16]), 
          .D1(n3242_adj_603), .CIN(n31060), .COUT(n31061), .S0(n3392_adj_2177[15]), 
          .S1(n3392_adj_2177[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_15.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_15.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_15.INJECT1_0 = "NO";
    defparam div_13_add_2249_15.INJECT1_1 = "NO";
    LUT4 rem_10_i1449_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[29]), 
         .D(n2140_adj_1790), .Z(n2239_adj_1832)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1449_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1455_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[23]), 
         .D(n2146_adj_1804), .Z(n2245_adj_1844)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1455_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_13 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[13]), 
          .D0(n3245_adj_720), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[14]), 
          .D1(n3244_adj_807), .CIN(n31059), .COUT(n31060), .S0(n3392_adj_2177[13]), 
          .S1(n3392_adj_2177[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_13.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_13.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_13.INJECT1_0 = "NO";
    defparam div_13_add_2249_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1458_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[20]), 
         .D(n2149_adj_1807), .Z(n2248_adj_1853)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1458_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1448_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[30]), 
         .D(n2139_adj_1785), .Z(n2238_adj_1833)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1448_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1457_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[21]), 
         .D(n2148_adj_1808), .Z(n2247_adj_1848)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1457_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1452_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[26]), 
         .D(n2143_adj_1793), .Z(n2242_adj_1841)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1452_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_11 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[11]), 
          .D0(n3247_adj_811), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[12]), 
          .D1(n3246_adj_736), .CIN(n31058), .COUT(n31059), .S0(n3392_adj_2177[11]), 
          .S1(n3392_adj_2177[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_11.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_11.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_11.INJECT1_0 = "NO";
    defparam div_13_add_2249_11.INJECT1_1 = "NO";
    LUT4 rem_10_i1454_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[24]), 
         .D(n2145_adj_1797), .Z(n2244_adj_1845)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1454_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_9 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[9]), 
          .D0(n3249_adj_698), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[10]), 
          .D1(n3248_adj_695), .CIN(n31057), .COUT(n31058), .S0(n3392_adj_2177[9]), 
          .S1(n3392_adj_2177[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_9.INIT0 = 16'hf1e0;
    defparam div_13_add_2249_9.INIT1 = 16'hf1e0;
    defparam div_13_add_2249_9.INJECT1_0 = "NO";
    defparam div_13_add_2249_9.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_7 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[7]), 
          .D0(n3251_adj_672), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[8]), 
          .D1(n3250_adj_704), .CIN(n31056), .COUT(n31057), .S0(n3392_adj_2177[7]), 
          .S1(n3392_adj_2177[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_7.INIT0 = 16'h0e1f;
    defparam div_13_add_2249_7.INIT1 = 16'hf1e0;
    defparam div_13_add_2249_7.INJECT1_0 = "NO";
    defparam div_13_add_2249_7.INJECT1_1 = "NO";
    LUT4 rem_10_i1463_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[15]), 
         .D(n2154_adj_1823), .Z(n2253_adj_1872)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1463_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_356 (.A(distance[8]), .B(distance[6]), .C(distance[11]), 
         .D(distance[9]), .Z(n34944)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_356.init = 16'hfffe;
    LUT4 div_9_i2187_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[28]), 
         .D(n3230), .Z(n3329_adj_2023)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2187_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2249_5 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[5]), 
          .D0(n3253_adj_657), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[6]), 
          .D1(n3252_adj_718), .CIN(n31055), .COUT(n31056), .S0(n3392_adj_2177[5]), 
          .S1(n3392_adj_2177[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_5.INIT0 = 16'hf1e0;
    defparam div_13_add_2249_5.INIT1 = 16'hf1e0;
    defparam div_13_add_2249_5.INJECT1_0 = "NO";
    defparam div_13_add_2249_5.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_3 (.A0(n13610), .B0(n28528), .C0(n3293_adj_2164[3]), 
          .D0(n348_adj_1735), .A1(n13610), .B1(n28528), .C1(n3293_adj_2164[4]), 
          .D1(n3254_adj_668), .CIN(n31054), .COUT(n31055), .S0(n3392_adj_2177[3]), 
          .S1(n3392_adj_2177[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_3.INIT0 = 16'hf1e0;
    defparam div_13_add_2249_3.INIT1 = 16'h0e1f;
    defparam div_13_add_2249_3.INJECT1_0 = "NO";
    defparam div_13_add_2249_3.INJECT1_1 = "NO";
    CCU2C div_13_add_2249_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n349), .B1(GND_net), .C1(GND_net), .D1(VCC_net), 
          .COUT(n31054), .S1(n3392_adj_2177[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2249_1.INIT0 = 16'h0000;
    defparam div_13_add_2249_1.INIT1 = 16'h555a;
    defparam div_13_add_2249_1.INJECT1_0 = "NO";
    defparam div_13_add_2249_1.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_29 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[30]), 
          .D0(n38192), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[31]), 
          .D1(n3128), .CIN(n31052), .S0(n3293_adj_2164[30]), .S1(n3293_adj_2164[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_29.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_29.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_29.INJECT1_0 = "NO";
    defparam div_13_add_2182_29.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_27 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[28]), 
          .D0(n3131), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[29]), 
          .D1(n38193), .CIN(n31051), .COUT(n31052), .S0(n3293_adj_2164[28]), 
          .S1(n3293_adj_2164[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_27.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_27.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_27.INJECT1_0 = "NO";
    defparam div_13_add_2182_27.INJECT1_1 = "NO";
    LUT4 div_9_i2067_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[14]), 
         .D(n3046), .Z(n3145)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2067_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2071_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[10]), 
         .D(n3050), .Z(n3149)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2071_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1464_3_lut_4_lut (.A(n28387), .B(n13597), .C(n2204_adj_2172[14]), 
         .D(n586), .Z(n2254_adj_1889)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1464_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2182_25 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[26]), 
          .D0(n3133), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[27]), 
          .D1(n38194), .CIN(n31050), .COUT(n31051), .S0(n3293_adj_2164[26]), 
          .S1(n3293_adj_2164[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_25.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_25.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_25.INJECT1_0 = "NO";
    defparam div_13_add_2182_25.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_23 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[24]), 
          .D0(n3135_adj_687), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[25]), 
          .D1(n3134_adj_794), .CIN(n31049), .COUT(n31050), .S0(n3293_adj_2164[24]), 
          .S1(n3293_adj_2164[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_23.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_23.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_23.INJECT1_0 = "NO";
    defparam div_13_add_2182_23.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_21 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[22]), 
          .D0(n3137_adj_674), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[23]), 
          .D1(n3136_adj_791), .CIN(n31048), .COUT(n31049), .S0(n3293_adj_2164[22]), 
          .S1(n3293_adj_2164[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_21.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_21.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_21.INJECT1_0 = "NO";
    defparam div_13_add_2182_21.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_19 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[20]), 
          .D0(n3139_adj_753), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[21]), 
          .D1(n3138_adj_661), .CIN(n31047), .COUT(n31048), .S0(n3293_adj_2164[20]), 
          .S1(n3293_adj_2164[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_19.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_19.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_19.INJECT1_0 = "NO";
    defparam div_13_add_2182_19.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_267 (.A(n28440), .B(n13590), .Z(n38272)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_rep_267.init = 16'heeee;
    LUT4 div_9_i1456_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[22]), 
         .D(n2147), .Z(n2246_adj_2018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1456_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1447_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[31]), 
         .D(n38274), .Z(n2237_adj_1916)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1447_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1462_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[16]), 
         .D(n2153), .Z(n2252_adj_2091)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1462_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1455_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[23]), 
         .D(n2146), .Z(n2245_adj_2015)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1455_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2182_17 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[18]), 
          .D0(n3141_adj_730), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[19]), 
          .D1(n3140_adj_772), .CIN(n31046), .COUT(n31047), .S0(n3293_adj_2164[18]), 
          .S1(n3293_adj_2164[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_17.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_17.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_17.INJECT1_0 = "NO";
    defparam div_13_add_2182_17.INJECT1_1 = "NO";
    LUT4 div_9_i1450_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[28]), 
         .D(n2141), .Z(n2240_adj_1922)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1450_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2182_15 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[16]), 
          .D0(n3143), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[17]), 
          .D1(n3142_adj_684), .CIN(n31045), .COUT(n31046), .S0(n3293_adj_2164[16]), 
          .S1(n3293_adj_2164[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_15.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_15.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_15.INJECT1_0 = "NO";
    defparam div_13_add_2182_15.INJECT1_1 = "NO";
    LUT4 div_9_i1451_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[27]), 
         .D(n2142), .Z(n2241_adj_1921)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1451_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1463_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[15]), 
         .D(n2154), .Z(n2253_adj_2092)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1463_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1452_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[26]), 
         .D(n2143), .Z(n2242_adj_1925)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1452_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1461_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[17]), 
         .D(n38278), .Z(n2251_adj_2089)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1461_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1449_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[29]), 
         .D(n2140), .Z(n2239_adj_1917)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1449_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1458_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[20]), 
         .D(n2149), .Z(n2248_adj_2086)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1458_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1459_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[19]), 
         .D(n2150), .Z(n2249_adj_2087)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1459_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1457_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[21]), 
         .D(n2148), .Z(n2247_adj_2017)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1457_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1460_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[18]), 
         .D(n2151), .Z(n2250_adj_2090)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1460_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2182_13 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[14]), 
          .D0(n3145_adj_806), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[15]), 
          .D1(n3144_adj_691), .CIN(n31044), .COUT(n31045), .S0(n3293_adj_2164[14]), 
          .S1(n3293_adj_2164[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_13.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_13.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_13.INJECT1_0 = "NO";
    defparam div_13_add_2182_13.INJECT1_1 = "NO";
    LUT4 div_9_i1453_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[25]), 
         .D(n2144), .Z(n2243_adj_1924)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1453_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1448_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[30]), 
         .D(n38275), .Z(n2238_adj_1918)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1448_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2182_11 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[12]), 
          .D0(n3147_adj_770), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[13]), 
          .D1(n3146_adj_768), .CIN(n31043), .COUT(n31044), .S0(n3293_adj_2164[12]), 
          .S1(n3293_adj_2164[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_11.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_11.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_11.INJECT1_0 = "NO";
    defparam div_13_add_2182_11.INJECT1_1 = "NO";
    LUT4 div_9_i2072_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[9]), 
         .D(n3051), .Z(n3150)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2072_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1454_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[24]), 
         .D(n38277), .Z(n2244_adj_2016)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1454_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1464_3_lut_4_lut (.A(n28440), .B(n13590), .C(n2204[14]), 
         .D(n337), .Z(n2254_adj_2093)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1464_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i14_3_lut (.A(n102), .B(n38[13]), .C(n3556), .Z(n338_adj_913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i14_3_lut.init = 16'hcaca;
    LUT4 div_9_i2060_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[21]), 
         .D(n3039), .Z(n3138)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2060_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i13_3_lut (.A(n105), .B(n38[12]), .C(n3556), .Z(n339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i13_3_lut.init = 16'hcaca;
    LUT4 div_9_i2063_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[18]), 
         .D(n3042), .Z(n3141)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2063_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_357 (.A(n1940_adj_1120), .B(n2006_adj_2182[31]), 
         .C(n38276), .D(n2041_adj_1109), .Z(n35714)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_357.init = 16'hffca;
    CCU2C div_13_add_2182_9 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[10]), 
          .D0(n3149_adj_694), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[11]), 
          .D1(n3148_adj_810), .CIN(n31042), .COUT(n31043), .S0(n3293_adj_2164[10]), 
          .S1(n3293_adj_2164[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_9.INIT0 = 16'hf1e0;
    defparam div_13_add_2182_9.INIT1 = 16'hf1e0;
    defparam div_13_add_2182_9.INJECT1_0 = "NO";
    defparam div_13_add_2182_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_358 (.A(n2039), .B(n2105[31]), .C(n38279), 
         .D(n2140), .Z(n36314)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_358.init = 16'hffca;
    LUT4 div_9_i2054_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[27]), 
         .D(n3033), .Z(n3132_adj_1728)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2054_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2182_7 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[8]), 
          .D0(n3151), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[9]), 
          .D1(n3150_adj_697), .CIN(n31041), .COUT(n31042), .S0(n3293_adj_2164[8]), 
          .S1(n3293_adj_2164[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_7.INIT0 = 16'h0e1f;
    defparam div_13_add_2182_7.INIT1 = 16'hf1e0;
    defparam div_13_add_2182_7.INJECT1_0 = "NO";
    defparam div_13_add_2182_7.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_5 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[6]), 
          .D0(n3153_adj_717), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[7]), 
          .D1(n3152_adj_671), .CIN(n31040), .COUT(n31041), .S0(n3293_adj_2164[6]), 
          .S1(n3293_adj_2164[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_5.INIT0 = 16'hf1e0;
    defparam div_13_add_2182_5.INIT1 = 16'hf1e0;
    defparam div_13_add_2182_5.INJECT1_0 = "NO";
    defparam div_13_add_2182_5.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_3 (.A0(n13614), .B0(n28522), .C0(n3194_adj_2167[4]), 
          .D0(n347_adj_667), .A1(n13614), .B1(n28522), .C1(n3194_adj_2167[5]), 
          .D1(n3154_adj_656), .CIN(n31039), .COUT(n31040), .S0(n3293_adj_2164[4]), 
          .S1(n3293_adj_2164[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_3.INIT0 = 16'hf1e0;
    defparam div_13_add_2182_3.INIT1 = 16'h0e1f;
    defparam div_13_add_2182_3.INJECT1_0 = "NO";
    defparam div_13_add_2182_3.INJECT1_1 = "NO";
    CCU2C div_13_add_2182_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n348_adj_1735), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n31039), .S1(n3293_adj_2164[3]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2182_1.INIT0 = 16'h0000;
    defparam div_13_add_2182_1.INIT1 = 16'h555a;
    defparam div_13_add_2182_1.INJECT1_0 = "NO";
    defparam div_13_add_2182_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_359 (.A(n2040), .B(n2105[30]), .C(n38279), 
         .D(n2141), .Z(n36310)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_359.init = 16'hffca;
    LUT4 i1_2_lut_rep_271 (.A(n28389), .B(n13636), .Z(n38276)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_rep_271.init = 16'heeee;
    LUT4 div_9_i2058_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[23]), 
         .D(n3037), .Z(n3136)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2058_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1313_3_lut_rep_268_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[31]), 
         .D(n1940_adj_1120), .Z(n38273)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1313_3_lut_rep_268_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1319_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[25]), 
         .D(n1946_adj_1128), .Z(n2045_adj_1048)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1319_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2064_3_lut_4_lut (.A(n28578), .B(n13548), .C(n3095[17]), 
         .D(n3043), .Z(n3142)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2064_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1316_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[28]), 
         .D(n1943_adj_1127), .Z(n2042_adj_1053)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1316_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_360 (.A(n3053_adj_1679), .B(n3095_adj_2184[7]), 
         .C(n38207), .D(n3151_adj_1294), .Z(n34812)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_360.init = 16'hca00;
    LUT4 div_13_i1321_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[23]), 
         .D(n1948_adj_1132), .Z(n2047_adj_1059)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1321_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1325_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[19]), 
         .D(n1952_adj_1145), .Z(n2051_adj_1061)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1325_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1317_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[27]), 
         .D(n1944_adj_1125), .Z(n2043_adj_1049)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1317_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_29 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[31]), 
          .D0(n3029_adj_1316), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n31038), .S0(n3194_adj_2167[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_29.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_29.INIT1 = 16'h0000;
    defparam div_13_add_2115_29.INJECT1_0 = "NO";
    defparam div_13_add_2115_29.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_27 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[29]), 
          .D0(n3031), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[30]), 
          .D1(n3030), .CIN(n31037), .COUT(n31038), .S0(n3194_adj_2167[29]), 
          .S1(n3194_adj_2167[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_27.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_27.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_27.INJECT1_0 = "NO";
    defparam div_13_add_2115_27.INJECT1_1 = "NO";
    LUT4 div_13_i1314_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[30]), 
         .D(n1941_adj_1126), .Z(n2040_adj_1051)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1314_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_361 (.A(n3036_adj_1673), .B(n3095_adj_2184[24]), 
         .C(n38207), .D(n3130_adj_2025), .Z(n35176)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_361.init = 16'hffca;
    LUT4 div_13_i1328_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[16]), 
         .D(n335_adj_1150), .Z(n2054_adj_1066)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1328_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1326_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[18]), 
         .D(n1953_adj_1151), .Z(n2052_adj_1063)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1326_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1327_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[17]), 
         .D(n1954_adj_1152), .Z(n2053_adj_1065)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1327_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24494_2_lut_rep_202 (.A(n28281), .B(n13628), .Z(n38207)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24494_2_lut_rep_202.init = 16'heeee;
    LUT4 div_13_i1323_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[21]), 
         .D(n1950_adj_1144), .Z(n2049_adj_1060)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1323_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_25 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[27]), 
          .D0(n3033_adj_1055), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[28]), 
          .D1(n3032_adj_1417), .CIN(n31036), .COUT(n31037), .S0(n3194_adj_2167[27]), 
          .S1(n3194_adj_2167[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_25.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_25.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_25.INJECT1_0 = "NO";
    defparam div_13_add_2115_25.INJECT1_1 = "NO";
    LUT4 rem_10_i2074_3_lut_rep_200_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[7]), 
         .D(n3053_adj_1679), .Z(n38205)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2074_3_lut_rep_200_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1320_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[24]), 
         .D(n1947_adj_1133), .Z(n2046_adj_1052)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1320_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2057_3_lut_rep_201_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[24]), 
         .D(n3036_adj_1673), .Z(n38206)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2057_3_lut_rep_201_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1322_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[22]), 
         .D(n1949_adj_1134), .Z(n2048_adj_1058)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1322_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2063_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[18]), 
         .D(n3042_adj_1653), .Z(n3141_adj_2075)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2063_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2050_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[31]), 
         .D(n38210), .Z(n3128_adj_2042)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2050_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1315_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[29]), 
         .D(n1942_adj_1121), .Z(n2041_adj_1109)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1315_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i20_3_lut (.A(n84), .B(n38[19]), .C(n3556), .Z(n332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i20_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2066_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[15]), 
         .D(n3045_adj_1633), .Z(n3144_adj_2067)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2066_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2053_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[28]), 
         .D(n3032_adj_1642), .Z(n3131_adj_2047)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2053_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2054_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[27]), 
         .D(n3033_adj_1670), .Z(n3132)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2054_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1318_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[26]), 
         .D(n1945_adj_1119), .Z(n2044_adj_1050)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1318_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_23 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[25]), 
          .D0(n3035_adj_1469), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[26]), 
          .D1(n38203), .CIN(n31035), .COUT(n31036), .S0(n3194_adj_2167[25]), 
          .S1(n3194_adj_2167[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_23.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_23.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_23.INJECT1_0 = "NO";
    defparam div_13_add_2115_23.INJECT1_1 = "NO";
    LUT4 div_13_i1324_3_lut_4_lut (.A(n28389), .B(n13636), .C(n2006_adj_2182[20]), 
         .D(n1951_adj_1143), .Z(n2050_adj_1062)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1324_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i76_3_lut (.A(n14790), .B(n197[0]), .C(n89[0]), .Z(duty2_14__N_473[0])) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(29[19:24])
    defparam i76_3_lut.init = 16'ha8a8;
    LUT4 i1_2_lut_4_lut_adj_362 (.A(n38281), .B(n2105[24]), .C(n38279), 
         .D(n2143), .Z(n36316)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_362.init = 16'hffca;
    LUT4 rem_10_i2061_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[20]), 
         .D(n3040_adj_1645), .Z(n3139_adj_2080)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2061_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1389_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[22]), 
         .D(n2048_adj_924), .Z(n2147_adj_1803)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1389_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1395_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[16]), 
         .D(n2054_adj_932), .Z(n2153_adj_1819)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1395_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_363 (.A(n35082), .B(n35068), .C(n2636), .D(n2646), 
         .Z(n13624)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_363.init = 16'hfffe;
    LUT4 i1_4_lut_adj_364 (.A(n2642), .B(n35078), .C(n35074), .D(n2637), 
         .Z(n35082)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_364.init = 16'hfffe;
    LUT4 i1_4_lut_adj_365 (.A(n2635), .B(n2644), .C(n2643), .D(n2645), 
         .Z(n35068)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_365.init = 16'hfffe;
    LUT4 i1_4_lut_adj_366 (.A(n2641), .B(n2640), .C(n2639), .D(n2638), 
         .Z(n35078)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_4_lut_adj_366.init = 16'hfffe;
    LUT4 i1_4_lut_adj_367 (.A(n2648), .B(n28293), .C(n2647), .D(n2649), 
         .Z(n28462)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_367.init = 16'h8000;
    LUT4 i24340_4_lut (.A(n2651), .B(n2650), .C(n28042), .D(n2652), 
         .Z(n28293)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i24340_4_lut.init = 16'heccc;
    LUT4 i24092_3_lut (.A(n342), .B(n2653), .C(n2654), .Z(n28042)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i24092_3_lut.init = 16'hecec;
    LUT4 div_9_i2197_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[18]), 
         .D(n3240), .Z(n3339_adj_875)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2197_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2060_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[21]), 
         .D(n3039_adj_1663), .Z(n3138_adj_2031)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2060_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1380_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[31]), 
         .D(n2039_adj_845), .Z(n2138_adj_1786)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1380_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1392_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[19]), 
         .D(n2051_adj_926), .Z(n2150_adj_1816)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1392_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1382_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[29]), 
         .D(n2041_adj_850), .Z(n2140_adj_1790)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1382_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2058_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[23]), 
         .D(n3037_adj_1667), .Z(n3136_adj_2097)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2058_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_21 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[23]), 
          .D0(n3037_adj_1475), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[24]), 
          .D1(n3036_adj_1176), .CIN(n31034), .COUT(n31035), .S0(n3194_adj_2167[23]), 
          .S1(n3194_adj_2167[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_21.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_21.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_21.INJECT1_0 = "NO";
    defparam div_13_add_2115_21.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_19 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[21]), 
          .D0(n3039_adj_1358), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[22]), 
          .D1(n3038_adj_1227), .CIN(n31033), .COUT(n31034), .S0(n3194_adj_2167[21]), 
          .S1(n3194_adj_2167[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_19.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_19.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_19.INJECT1_0 = "NO";
    defparam div_13_add_2115_19.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_17 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[19]), 
          .D0(n38208), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[20]), 
          .D1(n3040_adj_1116), .CIN(n31032), .COUT(n31033), .S0(n3194_adj_2167[19]), 
          .S1(n3194_adj_2167[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_17.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_17.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_17.INJECT1_0 = "NO";
    defparam div_13_add_2115_17.INJECT1_1 = "NO";
    LUT4 rem_10_i2055_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[26]), 
         .D(n3034_adj_1677), .Z(n3133_adj_2028)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2055_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1394_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[17]), 
         .D(n2053_adj_931), .Z(n2152_adj_1820)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1394_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_mux_3_i15_3_lut (.A(n99), .B(n38[14]), .C(n3556), .Z(n337_adj_1001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i15_3_lut.init = 16'hcaca;
    LUT4 rem_10_i2056_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[25]), 
         .D(n3035_adj_1657), .Z(n3134_adj_2070)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2056_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1391_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[20]), 
         .D(n2050_adj_927), .Z(n2149_adj_1807)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1391_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1381_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[30]), 
         .D(n2040_adj_844), .Z(n2139_adj_1785)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1381_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1390_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[21]), 
         .D(n2049_adj_925), .Z(n2148_adj_1808)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1390_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1385_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[26]), 
         .D(n2044_adj_905), .Z(n2143_adj_1793)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1385_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1383_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[28]), 
         .D(n2042_adj_849), .Z(n2141_adj_1789)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1383_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1387_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[24]), 
         .D(n2046), .Z(n2145_adj_1797)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1387_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1384_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[27]), 
         .D(n38280), .Z(n2142_adj_1794)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1384_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1386_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[25]), 
         .D(n2045_adj_922), .Z(n2144_adj_1798)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1386_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1393_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[18]), 
         .D(n2052_adj_928), .Z(n2151_adj_1815)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1393_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1388_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[23]), 
         .D(n2047_adj_923), .Z(n2146_adj_1804)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1388_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2052_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[29]), 
         .D(n3031_adj_1629), .Z(n3130_adj_2025)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2052_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_15 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[17]), 
          .D0(n3043_adj_1354), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[18]), 
          .D1(n3042_adj_1299), .CIN(n31031), .COUT(n31032), .S0(n3194_adj_2167[17]), 
          .S1(n3194_adj_2167[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_15.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_15.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_15.INJECT1_0 = "NO";
    defparam div_13_add_2115_15.INJECT1_1 = "NO";
    LUT4 rem_10_i2051_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[30]), 
         .D(n3030_adj_1665), .Z(n3129_adj_2036)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2051_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i2194_3_lut_4_lut (.A(n28492), .B(n13629), .C(n3293[21]), 
         .D(n3237), .Z(n3336_adj_808)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_9_i2194_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1396_3_lut_4_lut (.A(n28407), .B(n13595), .C(n2105_adj_2168[15]), 
         .D(n585), .Z(n2154_adj_1823)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1396_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2064_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[17]), 
         .D(n3043_adj_1639), .Z(n3142_adj_2101)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2064_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_368 (.A(n2053), .B(n2105[17]), .C(n38279), 
         .D(n2151), .Z(n35784)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_368.init = 16'hca00;
    LUT4 i1_2_lut_rep_274 (.A(n28263), .B(n13605), .Z(n38279)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_rep_274.init = 16'heeee;
    LUT4 div_9_i1394_3_lut_rep_273_4_lut (.A(n28263), .B(n13605), .C(n2105[17]), 
         .D(n2053), .Z(n38278)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1394_3_lut_rep_273_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1387_3_lut_rep_272_4_lut (.A(n28263), .B(n13605), .C(n2105[24]), 
         .D(n38281), .Z(n38277)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1387_3_lut_rep_272_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1381_3_lut_rep_270_4_lut (.A(n28263), .B(n13605), .C(n2105[30]), 
         .D(n2040), .Z(n38275)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1381_3_lut_rep_270_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1383_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[28]), 
         .D(n2042), .Z(n2141)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1383_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1393_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[18]), 
         .D(n2052), .Z(n2151)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1393_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_13 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[15]), 
          .D0(n3045_adj_1217), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[16]), 
          .D1(n3044_adj_1386), .CIN(n31030), .COUT(n31031), .S0(n3194_adj_2167[15]), 
          .S1(n3194_adj_2167[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_13.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_13.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_13.INJECT1_0 = "NO";
    defparam div_13_add_2115_13.INJECT1_1 = "NO";
    LUT4 div_13_mux_3_i12_3_lut (.A(n108), .B(n38[11]), .C(n3556), .Z(n340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_mux_3_i12_3_lut.init = 16'hcaca;
    CCU2C div_13_add_2115_11 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[13]), 
          .D0(n3047_adj_1398), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[14]), 
          .D1(n3046_adj_1449), .CIN(n31029), .COUT(n31030), .S0(n3194_adj_2167[13]), 
          .S1(n3194_adj_2167[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_11.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_11.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_11.INJECT1_0 = "NO";
    defparam div_13_add_2115_11.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_9 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[11]), 
          .D0(n3049_adj_1483), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[12]), 
          .D1(n3048_adj_1404), .CIN(n31028), .COUT(n31029), .S0(n3194_adj_2167[11]), 
          .S1(n3194_adj_2167[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_9.INIT0 = 16'hf1e0;
    defparam div_13_add_2115_9.INIT1 = 16'hf1e0;
    defparam div_13_add_2115_9.INJECT1_0 = "NO";
    defparam div_13_add_2115_9.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_7 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[9]), 
          .D0(n3051_adj_1382), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[10]), 
          .D1(n3050_adj_1181), .CIN(n31027), .COUT(n31028), .S0(n3194_adj_2167[9]), 
          .S1(n3194_adj_2167[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_7.INIT0 = 16'h0e1f;
    defparam div_13_add_2115_7.INIT1 = 16'hf1e0;
    defparam div_13_add_2115_7.INJECT1_0 = "NO";
    defparam div_13_add_2115_7.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_5 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[7]), 
          .D0(n3053_adj_1183), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[8]), 
          .D1(n3052_adj_1373), .CIN(n31026), .COUT(n31027), .S0(n3194_adj_2167[7]), 
          .S1(n3194_adj_2167[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_5.INIT0 = 16'hf1e0;
    defparam div_13_add_2115_5.INIT1 = 16'hf1e0;
    defparam div_13_add_2115_5.INJECT1_0 = "NO";
    defparam div_13_add_2115_5.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_369 (.A(n1842), .B(n35744), .C(n35746), .D(n1845), 
         .Z(n13600)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_369.init = 16'hfffe;
    LUT4 div_9_i1385_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[26]), 
         .D(n2044), .Z(n2143)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1385_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_370 (.A(n34766), .B(n34788), .C(n1850), .D(n27919), 
         .Z(n28359)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_370.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_371 (.A(n1847), .B(n1848), .C(n1849), .Z(n34766)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_371.init = 16'h8080;
    LUT4 rem_10_i2067_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[14]), 
         .D(n3046_adj_1651), .Z(n3145_adj_2040)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2067_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2062_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[19]), 
         .D(n3041_adj_1675), .Z(n3140_adj_2038)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2062_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23969_3_lut (.A(n583), .B(n1853), .C(n1854), .Z(n27919)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23969_3_lut.init = 16'hecec;
    LUT4 div_9_i1386_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[25]), 
         .D(n2045), .Z(n2144)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1386_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1380_3_lut_rep_269_4_lut (.A(n28263), .B(n13605), .C(n2105[31]), 
         .D(n2039), .Z(n38274)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1380_3_lut_rep_269_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2059_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[22]), 
         .D(n38215), .Z(n3137_adj_2096)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2059_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2076_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[5]), 
         .D(n595), .Z(n3154_adj_2106)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2076_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_372 (.A(n3), .B(n2[18]), .C(n27382), .D(n5), .Z(n582)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut_adj_372.init = 16'h4000;
    LUT4 div_9_i1388_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[23]), 
         .D(n2047), .Z(n2146)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1388_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1384_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[27]), 
         .D(n2043), .Z(n2142)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1384_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1391_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[20]), 
         .D(n2050), .Z(n2149)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1391_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_373 (.A(n27382), .B(n3), .C(n39), .Z(duty0_14__N_426[15])) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_adj_373.init = 16'h2020;
    LUT4 div_9_i1390_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[21]), 
         .D(n2049), .Z(n2148)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1390_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2115_3 (.A0(n13617), .B0(n28518), .C0(n3095_adj_2176[5]), 
          .D0(n346_adj_1140), .A1(n13617), .B1(n28518), .C1(n3095_adj_2176[6]), 
          .D1(n3054_adj_1265), .CIN(n31025), .COUT(n31026), .S0(n3194_adj_2167[5]), 
          .S1(n3194_adj_2167[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_3.INIT0 = 16'hf1e0;
    defparam div_13_add_2115_3.INIT1 = 16'h0e1f;
    defparam div_13_add_2115_3.INJECT1_0 = "NO";
    defparam div_13_add_2115_3.INJECT1_1 = "NO";
    CCU2C div_13_add_2115_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n347_adj_667), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n31025), .S1(n3194_adj_2167[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2115_1.INIT0 = 16'h0000;
    defparam div_13_add_2115_1.INIT1 = 16'h555a;
    defparam div_13_add_2115_1.INJECT1_0 = "NO";
    defparam div_13_add_2115_1.INJECT1_1 = "NO";
    PFUMX i62 (.BLUT(n60_adj_1030), .ALUT(n34594), .C0(n38307), .Z(n14790));
    PFUMX i16 (.BLUT(n34013), .ALUT(n34015), .C0(n38168), .Z(n5_adj_2103));
    PFUMX i62_adj_374 (.BLUT(n37_adj_1750), .ALUT(n34078), .C0(n38185), 
          .Z(n25_adj_2019));
    LUT4 div_9_i1389_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[22]), 
         .D(n2048), .Z(n2147)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1389_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i61 (.BLUT(n33434), .ALUT(n34474), .C0(n38197), .Z(n34));
    LUT4 div_9_i1396_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[15]), 
         .D(n336), .Z(n2154)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1396_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_27 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[30]), 
          .D0(n2931_adj_2115), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[31]), 
          .D1(n2930_adj_1583), .CIN(n31023), .S0(n3095_adj_2176[30]), 
          .S1(n3095_adj_2176[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_27.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_27.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_27.INJECT1_0 = "NO";
    defparam div_13_add_2048_27.INJECT1_1 = "NO";
    LUT4 rem_10_i2370_4_lut (.A(n3453), .B(n3568[3]), .C(n38307), .D(n3458), 
         .Z(n36[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2370_4_lut.init = 16'hc5ca;
    LUT4 rem_10_i2340_4_lut (.A(n3447), .B(n34936), .C(n3458), .D(n38175), 
         .Z(n3546)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B (C (D))))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2340_4_lut.init = 16'h6aaa;
    LUT4 div_9_i1382_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[29]), 
         .D(n2041), .Z(n2140)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1382_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2275_3_lut (.A(n3350), .B(n3392_adj_2163[7]), .C(n3359), 
         .Z(n3449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i2275_3_lut.init = 16'hcaca;
    L6MUX21 pwm_cnt_14__I_0_51_i30 (.D0(n24), .D1(n28), .SD(n36931), .Z(led_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    L6MUX21 pwm_cnt_14__I_0_52_i30 (.D0(n24_adj_609), .D1(n28_adj_1179), 
            .SD(n36874), .Z(led_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    L6MUX21 pwm_cnt_14__I_0_53_i30 (.D0(n24_adj_627), .D1(n28_adj_1407), 
            .SD(n36817), .Z(led_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    L6MUX21 pwm_cnt_14__I_0_54_i30 (.D0(n24_adj_654), .D1(n28_adj_1507), 
            .SD(n36760), .Z(led_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=4, LSE_RCOL=3, LSE_LLINE=370, LSE_RLINE=375 */ ;
    LUT4 div_9_i1392_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[19]), 
         .D(n2051), .Z(n2150)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1392_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_375 (.A(n3346), .B(n3338), .C(n3333), .D(n3337), 
         .Z(n34836)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_375.init = 16'hfffe;
    LUT4 div_13_i1257_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[20]), 
         .D(n1852_adj_1196), .Z(n1951_adj_1143)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1257_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1246_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[31]), 
         .D(n1841_adj_1187), .Z(n1940_adj_1120)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1246_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1395_3_lut_4_lut (.A(n28263), .B(n13605), .C(n2105[16]), 
         .D(n2054), .Z(n2153)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1395_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_376 (.A(n34872), .B(n598), .C(n3353), .D(n3354), 
         .Z(n33591)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_376.init = 16'ha8a0;
    LUT4 i1_4_lut_adj_377 (.A(n3234_adj_630), .B(n3229), .C(n3232_adj_1767), 
         .D(n3244_adj_551), .Z(n35286)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_377.init = 16'hfffe;
    LUT4 rem_10_i2071_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[10]), 
         .D(n3050_adj_1700), .Z(n3149_adj_2119)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2071_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1250_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[27]), 
         .D(n1845_adj_1379), .Z(n1944_adj_1125)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1250_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1260_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[17]), 
         .D(n334_adj_1199), .Z(n1954_adj_1152)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1260_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_25 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[28]), 
          .D0(n2933), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[29]), 
          .D1(n2932_adj_1546), .CIN(n31022), .COUT(n31023), .S0(n3095_adj_2176[28]), 
          .S1(n3095_adj_2176[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_25.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_25.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_25.INJECT1_0 = "NO";
    defparam div_13_add_2048_25.INJECT1_1 = "NO";
    CCU2C div_13_add_2048_23 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[26]), 
          .D0(n2935_adj_2114), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[27]), 
          .D1(n2934_adj_1556), .CIN(n31021), .COUT(n31022), .S0(n3095_adj_2176[26]), 
          .S1(n3095_adj_2176[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_23.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_23.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_23.INJECT1_0 = "NO";
    defparam div_13_add_2048_23.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_378 (.A(n34852), .B(n34710), .C(n33591), .D(n3350), 
         .Z(n3359)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i1_4_lut_adj_378.init = 16'heeea;
    LUT4 i1_4_lut_adj_379 (.A(n34836), .B(n34848), .C(n34846), .D(n34818), 
         .Z(n34852)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_379.init = 16'hfffe;
    LUT4 div_13_i1247_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[30]), 
         .D(n1842_adj_1190), .Z(n1941_adj_1126)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1247_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2075_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[6]), 
         .D(n3054_adj_1686), .Z(n3153_adj_2021)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2075_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_380 (.A(n34928), .B(n34812), .C(n3150_adj_2120), 
         .D(n27862), .Z(n28224)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_380.init = 16'ha8a0;
    LUT4 div_13_i1255_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[22]), 
         .D(n1850_adj_1195), .Z(n1949_adj_1134)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1255_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i2068_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[13]), 
         .D(n3047_adj_1690), .Z(n3146_adj_2073)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2068_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_381 (.A(n3147_adj_1996), .B(n3148_adj_2011), .C(n3149_adj_2119), 
         .Z(n34928)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_381.init = 16'h8080;
    LUT4 div_13_i1256_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[21]), 
         .D(n1851_adj_1194), .Z(n1950_adj_1144)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1256_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23913_3_lut (.A(n596), .B(n3153_adj_2021), .C(n3154_adj_2106), 
         .Z(n27862)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23913_3_lut.init = 16'hecec;
    LUT4 div_13_i1253_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[24]), 
         .D(n1848_adj_1191), .Z(n1947_adj_1133)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1253_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_382 (.A(n35192), .B(n35198), .C(n35188), .D(n35194), 
         .Z(n13619)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_382.init = 16'hfffe;
    LUT4 div_13_i1259_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[18]), 
         .D(n1854_adj_1201), .Z(n1953_adj_1151)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1259_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_383 (.A(n3146_adj_2073), .B(n3141_adj_2075), .C(n3131_adj_2047), 
         .D(n3143_adj_1297), .Z(n35192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_383.init = 16'hfffe;
    LUT4 i1_3_lut_adj_384 (.A(n3347), .B(n3348), .C(n3349), .Z(n34710)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_384.init = 16'h8080;
    LUT4 i1_4_lut_adj_385 (.A(n35176), .B(n35190), .C(n3132), .D(n3137_adj_2096), 
         .Z(n35198)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_385.init = 16'hfffe;
    LUT4 i1_3_lut_adj_386 (.A(n3138_adj_2031), .B(n3134_adj_2070), .C(n3129_adj_2036), 
         .Z(n35188)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_3_lut_adj_386.init = 16'hfefe;
    LUT4 rem_10_i2072_3_lut_4_lut (.A(n28281), .B(n13628), .C(n3095_adj_2184[9]), 
         .D(n3051_adj_1624), .Z(n3150_adj_2120)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam rem_10_i2072_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_387 (.A(n3133_adj_2028), .B(n3139_adj_2080), .C(n3128_adj_2042), 
         .D(n3144_adj_2067), .Z(n35194)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_387.init = 16'hfffe;
    LUT4 div_13_i1248_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[29]), 
         .D(n1843_adj_1189), .Z(n1942_adj_1121)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1248_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1249_3_lut_4_lut (.A(n28377), .B(n38283), .C(n1907_adj_2183[28]), 
         .D(n1844_adj_1188), .Z(n1943_adj_1127)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1249_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_388 (.A(n3140_adj_2038), .B(n3142_adj_2101), .C(n3136_adj_2097), 
         .D(n3145_adj_2040), .Z(n35190)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_388.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_389 (.A(n2942_adj_1592), .B(n2996_adj_2201[19]), 
         .C(n38209), .D(n3046_adj_1449), .Z(n35042)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_389.init = 16'hffca;
    LUT4 i24562_2_lut_rep_204 (.A(n28506), .B(n13618), .Z(n38209)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24562_2_lut_rep_204.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_390 (.A(n1947_adj_800), .B(n2006_adj_2170[24]), 
         .C(n38284), .D(n2040), .Z(n36046)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_390.init = 16'hffca;
    LUT4 div_13_i1995_3_lut_rep_203_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[19]), 
         .D(n2942_adj_1592), .Z(n38208)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1995_3_lut_rep_203_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_277 (.A(n28333), .B(n13604), .Z(n38282)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_rep_277.init = 16'heeee;
    LUT4 rem_10_i1317_3_lut_rep_275_4_lut (.A(n28333), .B(n13604), .C(n2006[27]), 
         .D(n1944), .Z(n38280)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1317_3_lut_rep_275_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1316_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[28]), 
         .D(n1943), .Z(n2042_adj_849)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1316_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1328_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[16]), 
         .D(n584), .Z(n2054_adj_932)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1328_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_391 (.A(n34700), .B(n34720), .C(n3050_adj_1700), 
         .D(n27878), .Z(n28281)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_391.init = 16'ha8a0;
    LUT4 rem_10_i1319_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[25]), 
         .D(n1946), .Z(n2045_adj_922)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1319_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_392 (.A(n3047_adj_1690), .B(n3048_adj_1692), .C(n3049_adj_1694), 
         .Z(n34700)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_392.init = 16'h8080;
    LUT4 i23929_3_lut (.A(n595), .B(n3053_adj_1679), .C(n3054_adj_1686), 
         .Z(n27878)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23929_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_393 (.A(n35162), .B(n35164), .C(n35156), .D(n35160), 
         .Z(n13628)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_393.init = 16'hfffe;
    CCU2C div_13_add_2048_21 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[24]), 
          .D0(n2937_adj_2113), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[25]), 
          .D1(n2936_adj_1577), .CIN(n31020), .COUT(n31021), .S0(n3095_adj_2176[24]), 
          .S1(n3095_adj_2176[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_21.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_21.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_21.INJECT1_0 = "NO";
    defparam div_13_add_2048_21.INJECT1_1 = "NO";
    CCU2C div_13_add_2048_19 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[22]), 
          .D0(n2939_adj_1579), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[23]), 
          .D1(n2938_adj_1618), .CIN(n31019), .COUT(n31020), .S0(n3095_adj_2176[22]), 
          .S1(n3095_adj_2176[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_19.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_19.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_19.INJECT1_0 = "NO";
    defparam div_13_add_2048_19.INJECT1_1 = "NO";
    CCU2C div_13_add_2048_17 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[20]), 
          .D0(n38213), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[21]), 
          .D1(n2940_adj_1501), .CIN(n31018), .COUT(n31019), .S0(n3095_adj_2176[20]), 
          .S1(n3095_adj_2176[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_17.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_17.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_17.INJECT1_0 = "NO";
    defparam div_13_add_2048_17.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_394 (.A(n3033_adj_1670), .B(n3036_adj_1673), .C(n3041_adj_1675), 
         .D(n3034_adj_1677), .Z(n35162)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_394.init = 16'hfffe;
    LUT4 div_13_i2005_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[9]), 
         .D(n2952_adj_2110), .Z(n3051_adj_1382)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2005_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_395 (.A(n3039_adj_1663), .B(n35142), .C(n35150), 
         .D(n3030_adj_1665), .Z(n35164)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_395.init = 16'hfffe;
    LUT4 rem_10_i1321_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[23]), 
         .D(n1948), .Z(n2047_adj_923)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1321_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_396 (.A(n3043_adj_1639), .B(n3037_adj_1667), .C(n3045_adj_1633), 
         .D(n3035_adj_1657), .Z(n35156)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_396.init = 16'hfffe;
    LUT4 i1_4_lut_adj_397 (.A(n3031_adj_1629), .B(n3042_adj_1653), .C(n3040_adj_1645), 
         .D(n3032_adj_1642), .Z(n35160)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_397.init = 16'hfffe;
    LUT4 rem_10_i1322_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[22]), 
         .D(n1949), .Z(n2048_adj_924)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1322_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_15 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[18]), 
          .D0(n2943_adj_1588), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[19]), 
          .D1(n2942_adj_1592), .CIN(n31017), .COUT(n31018), .S0(n3095_adj_2176[18]), 
          .S1(n3095_adj_2176[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_15.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_15.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_15.INJECT1_0 = "NO";
    defparam div_13_add_2048_15.INJECT1_1 = "NO";
    LUT4 div_13_i1992_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[22]), 
         .D(n2939_adj_1579), .Z(n3038_adj_1227)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1992_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1326_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[18]), 
         .D(n1953), .Z(n2052_adj_928)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1326_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1324_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[20]), 
         .D(n1951), .Z(n2050_adj_927)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1324_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_13 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[16]), 
          .D0(n2945_adj_1590), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[17]), 
          .D1(n2944_adj_2117), .CIN(n31016), .COUT(n31017), .S0(n3095_adj_2176[16]), 
          .S1(n3095_adj_2176[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_13.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_13.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_13.INJECT1_0 = "NO";
    defparam div_13_add_2048_13.INJECT1_1 = "NO";
    LUT4 rem_10_i1325_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[19]), 
         .D(n1952), .Z(n2051_adj_926)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1325_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1314_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[30]), 
         .D(n1941), .Z(n2040_adj_844)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1314_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1313_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[31]), 
         .D(n1940), .Z(n2039_adj_845)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1313_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_11 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[14]), 
          .D0(n2947_adj_1620), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[15]), 
          .D1(n2946_adj_2116), .CIN(n31015), .COUT(n31016), .S0(n3095_adj_2176[14]), 
          .S1(n3095_adj_2176[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_11.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_11.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_11.INJECT1_0 = "NO";
    defparam div_13_add_2048_11.INJECT1_1 = "NO";
    LUT4 div_13_i1999_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[15]), 
         .D(n2946_adj_2116), .Z(n3045_adj_1217)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1999_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1315_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[29]), 
         .D(n1942), .Z(n2041_adj_850)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1315_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_9 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[12]), 
          .D0(n2949_adj_1552), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[13]), 
          .D1(n2948_adj_1550), .CIN(n31014), .COUT(n31015), .S0(n3095_adj_2176[12]), 
          .S1(n3095_adj_2176[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_9.INIT0 = 16'hf1e0;
    defparam div_13_add_2048_9.INIT1 = 16'hf1e0;
    defparam div_13_add_2048_9.INJECT1_0 = "NO";
    defparam div_13_add_2048_9.INJECT1_1 = "NO";
    CCU2C div_13_add_2048_7 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[10]), 
          .D0(n2951_adj_1514), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[11]), 
          .D1(n2950_adj_1616), .CIN(n31013), .COUT(n31014), .S0(n3095_adj_2176[10]), 
          .S1(n3095_adj_2176[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_7.INIT0 = 16'h0e1f;
    defparam div_13_add_2048_7.INIT1 = 16'hf1e0;
    defparam div_13_add_2048_7.INJECT1_0 = "NO";
    defparam div_13_add_2048_7.INJECT1_1 = "NO";
    CCU2C div_13_add_2048_5 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[8]), 
          .D0(n2953_adj_1586), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[9]), 
          .D1(n2952_adj_2110), .CIN(n31012), .COUT(n31013), .S0(n3095_adj_2176[8]), 
          .S1(n3095_adj_2176[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_5.INIT0 = 16'hf1e0;
    defparam div_13_add_2048_5.INIT1 = 16'hf1e0;
    defparam div_13_add_2048_5.INJECT1_0 = "NO";
    defparam div_13_add_2048_5.INJECT1_1 = "NO";
    LUT4 div_13_i2007_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[7]), 
         .D(n2954_adj_2112), .Z(n3053_adj_1183)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2007_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_398 (.A(n34810), .B(n34692), .C(n2950), .D(n27888), 
         .Z(n28436)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_398.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_399 (.A(n2947_adj_571), .B(n2948), .C(n2949), .Z(n34810)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_399.init = 16'h8080;
    LUT4 div_13_i1984_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[30]), 
         .D(n2931_adj_2115), .Z(n3030)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1984_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23939_3_lut (.A(n594), .B(n2953), .C(n2954), .Z(n27888)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23939_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_400 (.A(n35226), .B(n35228), .C(n35220), .D(n35224), 
         .Z(n13592)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_400.init = 16'hfffe;
    LUT4 rem_10_i1327_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[17]), 
         .D(n1954), .Z(n2053_adj_931)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1327_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2006_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[8]), 
         .D(n2953_adj_1586), .Z(n3052_adj_1373)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2006_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_401 (.A(n2934), .B(n2930), .C(n2931_adj_535), .D(n2945), 
         .Z(n35226)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_401.init = 16'hfffe;
    LUT4 i1_4_lut_adj_402 (.A(n2942), .B(n35208), .C(n35206), .D(n2939), 
         .Z(n35228)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_402.init = 16'hfffe;
    LUT4 i1_3_lut_adj_403 (.A(n2932), .B(n2935), .C(n2944), .Z(n35220)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_3_lut_adj_403.init = 16'hfefe;
    LUT4 i1_4_lut_adj_404 (.A(n2943), .B(n2946), .C(n2936), .D(n2938), 
         .Z(n35224)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_404.init = 16'hfffe;
    LUT4 rem_10_i1323_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[21]), 
         .D(n1950), .Z(n2049_adj_925)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1323_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_2048_3 (.A0(n13618), .B0(n28506), .C0(n2996_adj_2201[6]), 
          .D0(n345_adj_2111), .A1(n13618), .B1(n28506), .C1(n2996_adj_2201[7]), 
          .D1(n2954_adj_2112), .CIN(n31011), .COUT(n31012), .S0(n3095_adj_2176[6]), 
          .S1(n3095_adj_2176[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_3.INIT0 = 16'hf1e0;
    defparam div_13_add_2048_3.INIT1 = 16'h0e1f;
    defparam div_13_add_2048_3.INJECT1_0 = "NO";
    defparam div_13_add_2048_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1318_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[26]), 
         .D(n1945), .Z(n2044_adj_905)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1318_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1987_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[27]), 
         .D(n2934_adj_1556), .Z(n3033_adj_1055)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1987_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1119_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[24]), 
         .D(n1353), .Z(n1749_adj_1436)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1119_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1320_3_lut_4_lut (.A(n28333), .B(n13604), .C(n2006[24]), 
         .D(n1947), .Z(n2046)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1320_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_405 (.A(n34658), .B(n34684), .C(n2850), .D(n27905), 
         .Z(n28307)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_405.init = 16'ha8a0;
    LUT4 i1_3_lut_rep_278 (.A(n35726), .B(n1846_adj_1384), .C(n1845_adj_1379), 
         .Z(n38283)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_3_lut_rep_278.init = 16'hfefe;
    LUT4 div_13_i1120_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[23]), 
         .D(n1354), .Z(n1750_adj_1443)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1120_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_279 (.A(n28526), .B(n13613), .Z(n38284)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_rep_279.init = 16'heeee;
    LUT4 div_13_i1988_3_lut_rep_198_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[26]), 
         .D(n2935_adj_2114), .Z(n38203)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1988_3_lut_rep_198_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1324_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[20]), 
         .D(n1951_adj_833), .Z(n2050)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1324_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1932_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[15]), 
         .D(n2847_adj_610), .Z(n2946_adj_2116)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1932_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_rep_284 (.A(n36346), .B(n1843), .C(n1845_adj_974), .Z(n38289)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_3_lut_rep_284.init = 16'hfefe;
    LUT4 div_9_i1327_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[17]), 
         .D(n1954_adj_863), .Z(n2053)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1327_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_adj_406 (.A(n2847), .B(n2848_adj_570), .C(n2849), .Z(n34658)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_406.init = 16'h8080;
    CCU2C div_13_add_2048_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n346_adj_1140), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n31011), .S1(n3095_adj_2176[5]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_2048_1.INIT0 = 16'h0000;
    defparam div_13_add_2048_1.INIT1 = 16'h555a;
    defparam div_13_add_2048_1.INJECT1_0 = "NO";
    defparam div_13_add_2048_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_280_4_lut (.A(n36346), .B(n1843), .C(n1845_adj_974), 
         .D(n28321), .Z(n38285)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_rep_280_4_lut.init = 16'hfffe;
    LUT4 div_13_i1921_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[26]), 
         .D(n2836_adj_628), .Z(n2935_adj_2114)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1921_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1990_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[24]), 
         .D(n2937_adj_2113), .Z(n3036_adj_1176)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1990_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23955_3_lut (.A(n593), .B(n2853), .C(n2854), .Z(n27905)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23955_3_lut.init = 16'hecec;
    LUT4 div_13_i2004_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[10]), 
         .D(n2951_adj_1514), .Z(n3050_adj_1181)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2004_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1313_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[31]), 
         .D(n1940_adj_758), .Z(n2039)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1313_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_407 (.A(n35440), .B(n35448), .C(n35424), .D(n35434), 
         .Z(n13598)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_407.init = 16'hfffe;
    LUT4 i1_4_lut_adj_408 (.A(n2843), .B(n2835), .C(n2832_adj_534), .D(n2842), 
         .Z(n35440)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_408.init = 16'hfffe;
    LUT4 div_9_i1321_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[23]), 
         .D(n1948_adj_829), .Z(n2047)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1321_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1325_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[19]), 
         .D(n1952_adj_840), .Z(n2051)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1325_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1317_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[27]), 
         .D(n1944_adj_785), .Z(n2043)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1317_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1938_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[9]), 
         .D(n2853_adj_591), .Z(n2952_adj_2110)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1938_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1917_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[30]), 
         .D(n2832_adj_592), .Z(n2931_adj_2115)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1917_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1985_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[29]), 
         .D(n2932_adj_1546), .Z(n3031)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1985_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1316_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[28]), 
         .D(n1943_adj_777), .Z(n2042)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1316_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_409 (.A(n35428), .B(n35444), .C(n2841), .D(n2838_adj_525), 
         .Z(n35448)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_409.init = 16'hfffe;
    CCU2C div_13_add_1981_27 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[31]), 
          .D0(n2831), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n31010), .S0(n2996_adj_2201[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_27.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_27.INIT1 = 16'h0000;
    defparam div_13_add_1981_27.INJECT1_0 = "NO";
    defparam div_13_add_1981_27.INJECT1_1 = "NO";
    CCU2C div_13_add_1981_25 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[29]), 
          .D0(n38219), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[30]), 
          .D1(n2832_adj_592), .CIN(n31009), .COUT(n31010), .S0(n2996_adj_2201[29]), 
          .S1(n2996_adj_2201[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_25.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_25.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_25.INJECT1_0 = "NO";
    defparam div_13_add_1981_25.INJECT1_1 = "NO";
    LUT4 div_9_i1319_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[25]), 
         .D(n1946_adj_802), .Z(n2045)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1319_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1320_3_lut_rep_276_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[24]), 
         .D(n1947_adj_800), .Z(n38281)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1320_3_lut_rep_276_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1996_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[18]), 
         .D(n2943_adj_1588), .Z(n3042_adj_1299)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1996_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1328_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[16]), 
         .D(n335), .Z(n2054)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1328_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_410 (.A(n2834), .B(n2845), .C(n2846), .D(n2833), 
         .Z(n35444)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_410.init = 16'hfffe;
    LUT4 div_9_i1322_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[22]), 
         .D(n1949_adj_827), .Z(n2048)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1322_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_411 (.A(n34728), .B(n34654), .C(n2750_adj_943), 
         .D(n27915), .Z(n28373)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_411.init = 16'ha8a0;
    LUT4 i1_3_lut_adj_412 (.A(n2747_adj_824), .B(n2748_adj_911), .C(n2749_adj_941), 
         .Z(n34728)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_412.init = 16'h8080;
    LUT4 div_9_i1315_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[29]), 
         .D(n1942_adj_779), .Z(n2041)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1315_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23965_3_lut (.A(n592), .B(n2753_adj_774), .C(n2754_adj_945), 
         .Z(n27915)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i23965_3_lut.init = 16'hecec;
    LUT4 i1_4_lut_adj_413 (.A(n35402), .B(n35420), .C(n35418), .D(n2741_adj_780), 
         .Z(n13626)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_413.init = 16'hfffe;
    LUT4 div_9_i1326_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[18]), 
         .D(n1953_adj_838), .Z(n2052)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1326_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1318_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[26]), 
         .D(n1945_adj_783), .Z(n2044)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1318_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1323_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[21]), 
         .D(n1950_adj_835), .Z(n2049)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1323_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_414 (.A(n2733_adj_884), .B(n35416), .C(n35410), 
         .D(n2735_adj_814), .Z(n35420)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_414.init = 16'hfffe;
    LUT4 i1_4_lut_adj_415 (.A(n2732_adj_648), .B(n2745), .C(n2743_adj_890), 
         .D(n2742_adj_892), .Z(n35418)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_415.init = 16'hfffe;
    LUT4 i1_4_lut_adj_416 (.A(n2740), .B(n2737_adj_798), .C(n2746_adj_818), 
         .D(n2738_adj_760), .Z(n35416)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_4_lut_adj_416.init = 16'hfffe;
    LUT4 div_9_i1314_3_lut_4_lut (.A(n28526), .B(n13613), .C(n2006_adj_2170[30]), 
         .D(n1941_adj_756), .Z(n2040)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1314_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1994_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[20]), 
         .D(n38213), .Z(n3040_adj_1116)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1994_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1180_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[30]), 
         .D(n1743_adj_1421), .Z(n1842_adj_1190)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1180_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1185_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[25]), 
         .D(n1748_adj_1438), .Z(n1847_adj_1192)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1185_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2001_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[13]), 
         .D(n2948_adj_1550), .Z(n3047_adj_1398)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2001_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1181_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[29]), 
         .D(n38286), .Z(n1843_adj_1189)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1181_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1187_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[23]), 
         .D(n1750_adj_1443), .Z(n1849_adj_1193)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1187_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1997_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[17]), 
         .D(n2944_adj_2117), .Z(n3043_adj_1354)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1997_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1191_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[19]), 
         .D(n1754_adj_1454), .Z(n1853_adj_1200)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1191_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1183_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[27]), 
         .D(n1746_adj_1432), .Z(n1845_adj_1379)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1183_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1192_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[18]), 
         .D(n333_adj_1452), .Z(n1854_adj_1201)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1192_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1993_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[21]), 
         .D(n2940_adj_1501), .Z(n3039_adj_1358)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1993_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i31818_2_lut_4_lut (.A(n38271), .B(n4540[12]), .C(n38307), .D(n89[9]), 
         .Z(n36650)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i31818_2_lut_4_lut.init = 16'hffca;
    LUT4 div_13_i1186_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[24]), 
         .D(n1749_adj_1436), .Z(n1848_adj_1191)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1186_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1981_23 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[27]), 
          .D0(n2835_adj_619), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[28]), 
          .D1(n2834_adj_640), .CIN(n31008), .COUT(n31009), .S0(n2996_adj_2201[27]), 
          .S1(n2996_adj_2201[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_23.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_23.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_23.INJECT1_0 = "NO";
    defparam div_13_add_1981_23.INJECT1_1 = "NO";
    CCU2C div_13_add_1981_21 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[25]), 
          .D0(n2837), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[26]), 
          .D1(n2836_adj_628), .CIN(n31007), .COUT(n31008), .S0(n2996_adj_2201[25]), 
          .S1(n2996_adj_2201[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_21.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_21.INJECT1_0 = "NO";
    defparam div_13_add_1981_21.INJECT1_1 = "NO";
    CCU2C div_13_add_1981_19 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[23]), 
          .D0(n2839_adj_643), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[24]), 
          .D1(n38222), .CIN(n31006), .COUT(n31007), .S0(n2996_adj_2201[23]), 
          .S1(n2996_adj_2201[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_19.INJECT1_0 = "NO";
    defparam div_13_add_1981_19.INJECT1_1 = "NO";
    LUT4 div_13_i1983_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[31]), 
         .D(n2930_adj_1583), .Z(n3029_adj_1316)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1983_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1188_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[22]), 
         .D(n1751_adj_1441), .Z(n1850_adj_1195)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1188_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1190_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[20]), 
         .D(n1753_adj_724), .Z(n1852_adj_1196)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1190_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_417 (.A(distance[15]), .B(distance[7]), .Z(n34942)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_417.init = 16'heeee;
    LUT4 div_13_i1179_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[31]), 
         .D(n1742_adj_1423), .Z(n1841_adj_1187)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1179_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1184_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[26]), 
         .D(n1747_adj_1430), .Z(n1846_adj_1384)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1184_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1189_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[21]), 
         .D(n38287), .Z(n1851_adj_1194)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1189_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1182_3_lut_4_lut (.A(n28566), .B(n13638), .C(n1808_adj_2185[28]), 
         .D(n1745_adj_1425), .Z(n1844_adj_1188)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1182_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i32317 (.BLUT(n37668), .ALUT(n37667), .C0(n38177), .Z(n37669));
    LUT4 div_9_i1259_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[18]), 
         .D(n1854_adj_968), .Z(n1953_adj_838)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1259_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1252_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[25]), 
         .D(n1847_adj_958), .Z(n1946_adj_802)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1252_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2008_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[6]), 
         .D(n345_adj_2111), .Z(n3054_adj_1265)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2008_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1251_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[26]), 
         .D(n1846_adj_956), .Z(n1945_adj_783)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1251_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1254_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[23]), 
         .D(n1849_adj_960), .Z(n1948_adj_829)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1254_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1250_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[27]), 
         .D(n1845_adj_974), .Z(n1944_adj_785)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1250_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1981_17 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[21]), 
          .D0(n2841_adj_616), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[22]), 
          .D1(n2840), .CIN(n31005), .COUT(n31006), .S0(n2996_adj_2201[21]), 
          .S1(n2996_adj_2201[22]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_17.INJECT1_0 = "NO";
    defparam div_13_add_1981_17.INJECT1_1 = "NO";
    LUT4 div_9_i1248_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[29]), 
         .D(n1843), .Z(n1942_adj_779)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1248_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1998_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[16]), 
         .D(n2945_adj_1590), .Z(n3044_adj_1386)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1998_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1981_15 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[19]), 
          .D0(n2843_adj_637), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[20]), 
          .D1(n2842_adj_620), .CIN(n31004), .COUT(n31005), .S0(n2996_adj_2201[19]), 
          .S1(n2996_adj_2201[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_15.INJECT1_0 = "NO";
    defparam div_13_add_1981_15.INJECT1_1 = "NO";
    CCU2C div_13_add_1981_13 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[17]), 
          .D0(n2845_adj_585), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[18]), 
          .D1(n38227), .CIN(n31003), .COUT(n31004), .S0(n2996_adj_2201[17]), 
          .S1(n2996_adj_2201[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_13.INJECT1_0 = "NO";
    defparam div_13_add_1981_13.INJECT1_1 = "NO";
    CCU2C div_13_add_1981_11 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[15]), 
          .D0(n2847_adj_610), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[16]), 
          .D1(n2846_adj_615), .CIN(n31002), .COUT(n31003), .S0(n2996_adj_2201[15]), 
          .S1(n2996_adj_2201[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_11.INJECT1_0 = "NO";
    defparam div_13_add_1981_11.INJECT1_1 = "NO";
    LUT4 div_9_i1256_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[21]), 
         .D(n1851_adj_963), .Z(n1950_adj_835)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1256_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1257_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[20]), 
         .D(n1852), .Z(n1951_adj_833)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1257_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2002_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[12]), 
         .D(n2949_adj_1552), .Z(n3048_adj_1404)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2002_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1260_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[17]), 
         .D(n334), .Z(n1954_adj_863)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1260_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1247_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[30]), 
         .D(n1842_adj_957), .Z(n1941_adj_756)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1247_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2413_3_lut_4_lut (.A(n28506), .B(n13618), .C(n3556), 
         .D(n4990[5]), .Z(n197[5])) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam div_13_i2413_3_lut_4_lut.init = 16'hfe0e;
    LUT4 div_13_i2000_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[14]), 
         .D(n2947_adj_1620), .Z(n3046_adj_1449)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2000_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1246_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[31]), 
         .D(n1841_adj_874), .Z(n1940_adj_758)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1246_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1258_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[19]), 
         .D(n1853_adj_967), .Z(n1952_adj_840)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1258_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1253_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[24]), 
         .D(n1848_adj_959), .Z(n1947_adj_800)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1253_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1249_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[28]), 
         .D(n1844), .Z(n1943_adj_777)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1249_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_9_i1255_3_lut_4_lut (.A(n28321), .B(n38289), .C(n1907_adj_2173[22]), 
         .D(n1850_adj_964), .Z(n1949_adj_827)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_i1255_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1981_9 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[13]), 
          .D0(n2849_adj_631), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[14]), 
          .D1(n2848_adj_646), .CIN(n31001), .COUT(n31002), .S0(n2996_adj_2201[13]), 
          .S1(n2996_adj_2201[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1981_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1981_9.INJECT1_0 = "NO";
    defparam div_13_add_1981_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1981_7 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[11]), 
          .D0(n2851_adj_647), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[12]), 
          .D1(n2850_adj_636), .CIN(n31000), .COUT(n31001), .S0(n2996_adj_2201[11]), 
          .S1(n2996_adj_2201[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1981_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1981_7.INJECT1_0 = "NO";
    defparam div_13_add_1981_7.INJECT1_1 = "NO";
    LUT4 rem_10_i1249_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[28]), 
         .D(n38291), .Z(n1943)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1249_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1986_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[28]), 
         .D(n2933), .Z(n3032_adj_1417)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1986_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1250_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[27]), 
         .D(n1845), .Z(n1944)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1250_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1991_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[23]), 
         .D(n2938_adj_1618), .Z(n3037_adj_1475)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1991_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i2003_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[11]), 
         .D(n2950_adj_1616), .Z(n3049_adj_1483)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i2003_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1255_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[22]), 
         .D(n1850), .Z(n1949)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1255_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1258_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[19]), 
         .D(n1853), .Z(n1952)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1258_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1246_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[31]), 
         .D(n1841), .Z(n1940)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1246_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1989_3_lut_4_lut (.A(n28506), .B(n13618), .C(n2996_adj_2201[25]), 
         .D(n2936_adj_1577), .Z(n3035_adj_1469)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1989_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1981_5 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[9]), 
          .D0(n2853_adj_591), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[10]), 
          .D1(n2852), .CIN(n30999), .COUT(n31000), .S0(n2996_adj_2201[9]), 
          .S1(n2996_adj_2201[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1981_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1981_5.INJECT1_0 = "NO";
    defparam div_13_add_1981_5.INJECT1_1 = "NO";
    LUT4 rem_10_i1248_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[29]), 
         .D(n38290), .Z(n1942)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1248_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1252_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[25]), 
         .D(n1847), .Z(n1946)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1252_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1259_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[18]), 
         .D(n1854), .Z(n1953)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1259_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1260_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[17]), 
         .D(n583), .Z(n1954)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1260_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_418 (.A(n2930), .B(n2996_adj_2193[31]), .C(n38217), 
         .D(n3046_adj_1651), .Z(n35150)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam i1_2_lut_4_lut_adj_418.init = 16'hffca;
    LUT4 rem_10_i1254_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[23]), 
         .D(n1849), .Z(n1948)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1254_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1257_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[20]), 
         .D(n38292), .Z(n1951)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1257_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1247_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[30]), 
         .D(n1842), .Z(n1941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1247_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_419 (.A(n2932_adj_709), .B(n2996[29]), .C(n38218), 
         .D(n3035), .Z(n35992)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_419.init = 16'hffca;
    CCU2C div_13_add_1981_3 (.A0(n13621), .B0(n28484), .C0(n2897_adj_2189[7]), 
          .D0(n344_adj_2118), .A1(n13621), .B1(n28484), .C1(n2897_adj_2189[8]), 
          .D1(n2854_adj_601), .CIN(n30998), .COUT(n30999), .S0(n2996_adj_2201[7]), 
          .S1(n2996_adj_2201[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1981_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1981_3.INJECT1_0 = "NO";
    defparam div_13_add_1981_3.INJECT1_1 = "NO";
    LUT4 rem_10_i1256_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[21]), 
         .D(n1851), .Z(n1950)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1256_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1251_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[26]), 
         .D(n1846), .Z(n1945)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1251_3_lut_4_lut.init = 16'hf1e0;
    LUT4 rem_10_i1253_3_lut_4_lut (.A(n28359), .B(n13600), .C(n1907[24]), 
         .D(n1848), .Z(n1947)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_i1253_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_420 (.A(distance[5]), .B(distance[4]), .Z(n34774)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_420.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_421 (.A(n1645), .B(n1709_adj_2169[29]), .C(n38288), 
         .D(n1743_adj_1421), .Z(n35728)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_421.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_422 (.A(n2931), .B(n2996[30]), .C(n38218), 
         .D(n3039), .Z(n35982)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam i1_2_lut_4_lut_adj_422.init = 16'hffca;
    LUT4 i1_2_lut_4_lut_adj_423 (.A(n2842_adj_620), .B(n2897_adj_2189[20]), 
         .C(n38214), .D(n2932_adj_1546), .Z(n35240)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_423.init = 16'hffca;
    PFUMX i32456 (.BLUT(n38058), .ALUT(n38057), .C0(n3359), .Z(n38059));
    LUT4 i1_2_lut_4_lut_adj_424 (.A(n330), .B(n1709_adj_2169[21]), .C(n38288), 
         .D(n1751_adj_1441), .Z(n34790)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_4_lut_adj_424.init = 16'hca00;
    LUT4 i1_2_lut_adj_425 (.A(distance[3]), .B(distance[2]), .Z(n34772)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_425.init = 16'heeee;
    LUT4 i1_2_lut_rep_283 (.A(n28562), .B(n13640), .Z(n38288)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam i1_2_lut_rep_283.init = 16'heeee;
    LUT4 div_13_i1122_3_lut_rep_282_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[21]), 
         .D(n330), .Z(n38287)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1122_3_lut_rep_282_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1114_3_lut_rep_281_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[29]), 
         .D(n1645), .Z(n38286)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1114_3_lut_rep_281_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_426 (.A(n38353), .B(n34129), .C(n38352), .D(n34970), 
         .Z(n3)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_426.init = 16'hfffe;
    CCU2C div_13_add_1981_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n345_adj_2111), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30998), .S1(n2996_adj_2201[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1981_1.INIT0 = 16'h0000;
    defparam div_13_add_1981_1.INIT1 = 16'h555a;
    defparam div_13_add_1981_1.INJECT1_0 = "NO";
    defparam div_13_add_1981_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_25 (.A0(n13622), .B0(n28468), .C0(n2798[30]), 
          .D0(n2733), .A1(n13622), .B1(n28468), .C1(n2798[31]), .D1(n2732), 
          .CIN(n30996), .S0(n2897_adj_2189[30]), .S1(n2897_adj_2189[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_25.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_25.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_25.INJECT1_0 = "NO";
    defparam div_13_add_1914_25.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_23 (.A0(n13622), .B0(n28468), .C0(n2798[28]), 
          .D0(n2735), .A1(n13622), .B1(n28468), .C1(n2798[29]), .D1(n2734), 
          .CIN(n30995), .COUT(n30996), .S0(n2897_adj_2189[28]), .S1(n2897_adj_2189[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_23.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_23.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_23.INJECT1_0 = "NO";
    defparam div_13_add_1914_23.INJECT1_1 = "NO";
    LUT4 i24544_2_lut_rep_209 (.A(n28484), .B(n13621), .Z(n38214)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i24544_2_lut_rep_209.init = 16'heeee;
    LUT4 div_13_i1115_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[28]), 
         .D(n1448), .Z(n1745_adj_1425)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1115_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1930_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[17]), 
         .D(n2845_adj_585), .Z(n2944_adj_2117)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1930_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_427 (.A(n34966), .B(n10_adj_2159), .C(distance[8]), 
         .D(distance[7]), .Z(n34129)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_427.init = 16'h8000;
    LUT4 div_13_i1118_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[25]), 
         .D(n1352), .Z(n1748_adj_1438)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1118_3_lut_4_lut.init = 16'hf1e0;
    LUT4 div_13_i1124_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[19]), 
         .D(n332), .Z(n1754_adj_1454)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1124_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i32260 (.BLUT(n37487), .ALUT(n37486), .C0(n38168), .Z(n37488));
    CCU2C add_1401_11 (.A0(n28331), .B0(n13553), .C0(GND_net), .D0(VCC_net), 
          .A1(n28319), .B1(n13554), .C1(GND_net), .D1(VCC_net), .CIN(n30819), 
          .COUT(n30820), .S0(n4540[9]), .S1(n4540[10]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_11.INIT0 = 16'h1111;
    defparam add_1401_11.INIT1 = 16'h1111;
    defparam add_1401_11.INJECT1_0 = "NO";
    defparam add_1401_11.INJECT1_1 = "NO";
    CCU2C rem_10_add_1244_13 (.A0(n13631), .B0(n28090), .C0(n1808[27]), 
          .D0(n1746), .A1(n13631), .B1(n28090), .C1(n1808[28]), .D1(n1745_adj_1502), 
          .CIN(n30609), .COUT(n30610), .S0(n1907[27]), .S1(n1907[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(70[20:34])
    defparam rem_10_add_1244_13.INIT0 = 16'h0e1f;
    defparam rem_10_add_1244_13.INIT1 = 16'h0e1f;
    defparam rem_10_add_1244_13.INJECT1_0 = "NO";
    defparam rem_10_add_1244_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_428 (.A(distance[15]), .B(distance[11]), .Z(n34970)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_428.init = 16'heeee;
    LUT4 div_13_i1940_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[7]), 
         .D(n344_adj_2118), .Z(n2954_adj_2112)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1940_3_lut_4_lut.init = 16'hf1e0;
    CCU2C add_1401_9 (.A0(n28554), .B0(n13551), .C0(GND_net), .D0(VCC_net), 
          .A1(n28544), .B1(n13552), .C1(GND_net), .D1(VCC_net), .CIN(n30818), 
          .COUT(n30819), .S0(n4540[7]), .S1(n4540[8]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_9.INIT0 = 16'h1111;
    defparam add_1401_9.INIT1 = 16'h1111;
    defparam add_1401_9.INJECT1_0 = "NO";
    defparam add_1401_9.INJECT1_1 = "NO";
    CCU2C add_1401_7 (.A0(n28574), .B0(n13549), .C0(GND_net), .D0(VCC_net), 
          .A1(n28568), .B1(n13550), .C1(GND_net), .D1(VCC_net), .CIN(n30817), 
          .COUT(n30818), .S0(n4540[5]), .S1(n4540[6]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_7.INIT0 = 16'h1111;
    defparam add_1401_7.INIT1 = 16'h1111;
    defparam add_1401_7.INJECT1_0 = "NO";
    defparam add_1401_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_21 (.A0(n13622), .B0(n28468), .C0(n2798[26]), 
          .D0(n2737), .A1(n13622), .B1(n28468), .C1(n2798[27]), .D1(n2736), 
          .CIN(n30994), .COUT(n30995), .S0(n2897_adj_2189[26]), .S1(n2897_adj_2189[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_21.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_21.INJECT1_0 = "NO";
    defparam div_13_add_1914_21.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_9 (.A0(n13557), .B0(n28269), .C0(n2303[19]), 
          .D0(n2249_adj_2087), .A1(n13557), .B1(n28269), .C1(n2303[20]), 
          .D1(n2248_adj_2086), .CIN(n30693), .COUT(n30694), .S0(n2402_adj_2195[19]), 
          .S1(n2402_adj_2195[20]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_9.INIT0 = 16'hf1e0;
    defparam div_9_add_1579_9.INIT1 = 16'hf1e0;
    defparam div_9_add_1579_9.INJECT1_0 = "NO";
    defparam div_9_add_1579_9.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_19 (.A0(n13622), .B0(n28468), .C0(n2798[24]), 
          .D0(n2739), .A1(n13622), .B1(n28468), .C1(n2798[25]), .D1(n2738), 
          .CIN(n30993), .COUT(n30994), .S0(n2897_adj_2189[24]), .S1(n2897_adj_2189[25]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_19.INJECT1_0 = "NO";
    defparam div_13_add_1914_19.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_7 (.A0(n13557), .B0(n28269), .C0(n2303[17]), 
          .D0(n2251_adj_2089), .A1(n13557), .B1(n28269), .C1(n2303[18]), 
          .D1(n2250_adj_2090), .CIN(n30692), .COUT(n30693), .S0(n2402_adj_2195[17]), 
          .S1(n2402_adj_2195[18]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_7.INIT0 = 16'h0e1f;
    defparam div_9_add_1579_7.INIT1 = 16'hf1e0;
    defparam div_9_add_1579_7.INJECT1_0 = "NO";
    defparam div_9_add_1579_7.INJECT1_1 = "NO";
    CCU2C add_1401_5 (.A0(n28588), .B0(n13547), .C0(GND_net), .D0(VCC_net), 
          .A1(n28578), .B1(n13548), .C1(GND_net), .D1(VCC_net), .CIN(n30816), 
          .COUT(n30817), .S0(n4540[3]), .S1(n4540[4]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_5.INIT0 = 16'h1111;
    defparam add_1401_5.INIT1 = 16'h1111;
    defparam add_1401_5.INJECT1_0 = "NO";
    defparam add_1401_5.INJECT1_1 = "NO";
    CCU2C add_1401_3 (.A0(n28512), .B0(n13602), .C0(GND_net), .D0(VCC_net), 
          .A1(n28492), .B1(n13629), .C1(GND_net), .D1(VCC_net), .CIN(n30815), 
          .COUT(n30816), .S0(n4540[1]), .S1(n4540[2]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_3.INIT0 = 16'h1111;
    defparam add_1401_3.INIT1 = 16'h1111;
    defparam add_1401_3.INJECT1_0 = "NO";
    defparam add_1401_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_17 (.A0(n13622), .B0(n28468), .C0(n2798[22]), 
          .D0(n2741), .A1(n13622), .B1(n28468), .C1(n2798[23]), .D1(n38233), 
          .CIN(n30992), .COUT(n30993), .S0(n2897_adj_2189[22]), .S1(n2897_adj_2189[23]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_17.INJECT1_0 = "NO";
    defparam div_13_add_1914_17.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_15 (.A0(n13622), .B0(n28468), .C0(n2798[20]), 
          .D0(n2743), .A1(n13622), .B1(n28468), .C1(n2798[21]), .D1(n2742), 
          .CIN(n30991), .COUT(n30992), .S0(n2897_adj_2189[20]), .S1(n2897_adj_2189[21]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_15.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_15.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_15.INJECT1_0 = "NO";
    defparam div_13_add_1914_15.INJECT1_1 = "NO";
    CCU2C add_1401_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(VCC_net), 
          .A1(n28160), .B1(n13556), .C1(GND_net), .D1(VCC_net), .COUT(n30815), 
          .S1(n4540[0]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam add_1401_1.INIT0 = 16'h0000;
    defparam add_1401_1.INIT1 = 16'heee1;
    defparam add_1401_1.INJECT1_0 = "NO";
    defparam add_1401_1.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_5 (.A0(n13557), .B0(n28269), .C0(n2303[15]), 
          .D0(n2253_adj_2092), .A1(n13557), .B1(n28269), .C1(n2303[16]), 
          .D1(n2252_adj_2091), .CIN(n30691), .COUT(n30692), .S0(n2402_adj_2195[15]), 
          .S1(n2402_adj_2195[16]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_5.INIT0 = 16'hf1e0;
    defparam div_9_add_1579_5.INIT1 = 16'hf1e0;
    defparam div_9_add_1579_5.INJECT1_0 = "NO";
    defparam div_9_add_1579_5.INJECT1_1 = "NO";
    CCU2C div_9_add_2182_29 (.A0(n13547), .B0(n28588), .C0(n3194[30]), 
          .D0(n3129), .A1(n13547), .B1(n28588), .C1(n3194[31]), .D1(n3128_adj_1528), 
          .CIN(n30813), .S0(n3293[30]), .S1(n3293[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_29.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_29.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_29.INJECT1_0 = "NO";
    defparam div_9_add_2182_29.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_13 (.A0(n13622), .B0(n28468), .C0(n2798[18]), 
          .D0(n38232), .A1(n13622), .B1(n28468), .C1(n2798[19]), .D1(n2744), 
          .CIN(n30990), .COUT(n30991), .S0(n2897_adj_2189[18]), .S1(n2897_adj_2189[19]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_13.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_13.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_13.INJECT1_0 = "NO";
    defparam div_13_add_1914_13.INJECT1_1 = "NO";
    PFUMX i32506 (.BLUT(n38416), .ALUT(n38417), .C0(n38307), .Z(n38418));
    CCU2C div_13_add_1914_11 (.A0(n13622), .B0(n28468), .C0(n2798[16]), 
          .D0(n2747), .A1(n13622), .B1(n28468), .C1(n2798[17]), .D1(n2746), 
          .CIN(n30989), .COUT(n30990), .S0(n2897_adj_2189[16]), .S1(n2897_adj_2189[17]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_11.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_11.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_11.INJECT1_0 = "NO";
    defparam div_13_add_1914_11.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_9 (.A0(n13622), .B0(n28468), .C0(n2798[14]), 
          .D0(n2749), .A1(n13622), .B1(n28468), .C1(n2798[15]), .D1(n2748), 
          .CIN(n30988), .COUT(n30989), .S0(n2897_adj_2189[14]), .S1(n2897_adj_2189[15]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_9.INIT0 = 16'hf1e0;
    defparam div_13_add_1914_9.INIT1 = 16'hf1e0;
    defparam div_13_add_1914_9.INJECT1_0 = "NO";
    defparam div_13_add_1914_9.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_429 (.A(distance[9]), .B(distance[6]), .C(distance[5]), 
         .Z(n34966)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_429.init = 16'h8080;
    CCU2C div_9_add_1579_3 (.A0(n13557), .B0(n28269), .C0(n2303[13]), 
          .D0(n338), .A1(n13557), .B1(n28269), .C1(n2303[14]), .D1(n2254_adj_2093), 
          .CIN(n30690), .COUT(n30691), .S0(n2402_adj_2195[13]), .S1(n2402_adj_2195[14]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_3.INIT0 = 16'hf1e0;
    defparam div_9_add_1579_3.INIT1 = 16'h0e1f;
    defparam div_9_add_1579_3.INJECT1_0 = "NO";
    defparam div_9_add_1579_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_7 (.A0(n13622), .B0(n28468), .C0(n2798[12]), 
          .D0(n2751), .A1(n13622), .B1(n28468), .C1(n2798[13]), .D1(n2750), 
          .CIN(n30987), .COUT(n30988), .S0(n2897_adj_2189[12]), .S1(n2897_adj_2189[13]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_7.INIT0 = 16'h0e1f;
    defparam div_13_add_1914_7.INIT1 = 16'hf1e0;
    defparam div_13_add_1914_7.INJECT1_0 = "NO";
    defparam div_13_add_1914_7.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_5 (.A0(n13622), .B0(n28468), .C0(n2798[10]), 
          .D0(n2753), .A1(n13622), .B1(n28468), .C1(n2798[11]), .D1(n2752), 
          .CIN(n30986), .COUT(n30987), .S0(n2897_adj_2189[10]), .S1(n2897_adj_2189[11]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_5.INIT0 = 16'hf1e0;
    defparam div_13_add_1914_5.INIT1 = 16'hf1e0;
    defparam div_13_add_1914_5.INJECT1_0 = "NO";
    defparam div_13_add_1914_5.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_3 (.A0(n13622), .B0(n28468), .C0(n2798[8]), 
          .D0(n343), .A1(n13622), .B1(n28468), .C1(n2798[9]), .D1(n2754), 
          .CIN(n30985), .COUT(n30986), .S0(n2897_adj_2189[8]), .S1(n2897_adj_2189[9]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_3.INIT0 = 16'hf1e0;
    defparam div_13_add_1914_3.INIT1 = 16'h0e1f;
    defparam div_13_add_1914_3.INJECT1_0 = "NO";
    defparam div_13_add_1914_3.INJECT1_1 = "NO";
    CCU2C div_13_add_1914_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n344_adj_2118), .B1(GND_net), .C1(GND_net), 
          .D1(VCC_net), .COUT(n30985), .S1(n2897_adj_2189[7]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1914_1.INIT0 = 16'h0000;
    defparam div_13_add_1914_1.INIT1 = 16'h555a;
    defparam div_13_add_1914_1.INJECT1_0 = "NO";
    defparam div_13_add_1914_1.INJECT1_1 = "NO";
    CCU2C div_13_add_1847_25 (.A0(n13624), .B0(n28462), .C0(n2699[31]), 
          .D0(n38241), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n30984), .S0(n2798[31]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_25.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_25.INIT1 = 16'h0000;
    defparam div_13_add_1847_25.INJECT1_0 = "NO";
    defparam div_13_add_1847_25.INJECT1_1 = "NO";
    CCU2C div_13_add_1847_23 (.A0(n13624), .B0(n28462), .C0(n2699[29]), 
          .D0(n2635), .A1(n13624), .B1(n28462), .C1(n2699[30]), .D1(n2634), 
          .CIN(n30983), .COUT(n30984), .S0(n2798[29]), .S1(n2798[30]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_23.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_23.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_23.INJECT1_0 = "NO";
    defparam div_13_add_1847_23.INJECT1_1 = "NO";
    PFUMX i32504 (.BLUT(n38413), .ALUT(n38414), .C0(n66_adj_2), .Z(n1352));
    CCU2C div_9_add_2182_27 (.A0(n13547), .B0(n28588), .C0(n3194[28]), 
          .D0(n3131_adj_1727), .A1(n13547), .B1(n28588), .C1(n3194[29]), 
          .D1(n3130), .CIN(n30812), .COUT(n30813), .S0(n3293[28]), .S1(n3293[29]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_27.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_27.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_27.INJECT1_0 = "NO";
    defparam div_9_add_2182_27.INJECT1_1 = "NO";
    LUT4 div_13_i1121_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[22]), 
         .D(n329), .Z(n1751_adj_1441)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1121_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1847_21 (.A0(n13624), .B0(n28462), .C0(n2699[27]), 
          .D0(n2637), .A1(n13624), .B1(n28462), .C1(n2699[28]), .D1(n2636), 
          .CIN(n30982), .COUT(n30983), .S0(n2798[27]), .S1(n2798[28]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_21.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_21.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_21.INJECT1_0 = "NO";
    defparam div_13_add_1847_21.INJECT1_1 = "NO";
    PFUMX i32265 (.BLUT(n37505), .ALUT(n37504), .C0(n38168), .Z(n37506));
    LUT4 div_13_i1116_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[27]), 
         .D(n1350), .Z(n1746_adj_1432)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1116_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1847_19 (.A0(n13624), .B0(n28462), .C0(n2699[25]), 
          .D0(n2639), .A1(n13624), .B1(n28462), .C1(n2699[26]), .D1(n2638), 
          .CIN(n30981), .COUT(n30982), .S0(n2798[25]), .S1(n2798[26]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_19.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_19.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_19.INJECT1_0 = "NO";
    defparam div_13_add_1847_19.INJECT1_1 = "NO";
    PFUMX i32502 (.BLUT(n38410), .ALUT(n38411), .C0(n69_adj_6), .Z(n1353));
    LUT4 i1183_2_lut (.A(distance[3]), .B(distance[4]), .Z(n10_adj_2159)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1183_2_lut.init = 16'heeee;
    CCU2C div_9_add_2182_25 (.A0(n13547), .B0(n28588), .C0(n3194[26]), 
          .D0(n3133_adj_2014), .A1(n13547), .B1(n28588), .C1(n3194[27]), 
          .D1(n3132_adj_1728), .CIN(n30811), .COUT(n30812), .S0(n3293[26]), 
          .S1(n3293[27]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_2182_25.INIT0 = 16'h0e1f;
    defparam div_9_add_2182_25.INIT1 = 16'h0e1f;
    defparam div_9_add_2182_25.INJECT1_0 = "NO";
    defparam div_9_add_2182_25.INJECT1_1 = "NO";
    CCU2C div_9_add_1579_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(VCC_net), .A1(n12154), .B1(n5), .C1(n54), .D1(n35[12]), 
          .COUT(n30690), .S1(n2402_adj_2195[12]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(69[15:29])
    defparam div_9_add_1579_1.INIT0 = 16'h0000;
    defparam div_9_add_1579_1.INIT1 = 16'habef;
    defparam div_9_add_1579_1.INJECT1_0 = "NO";
    defparam div_9_add_1579_1.INJECT1_1 = "NO";
    LUT4 div_13_i1923_3_lut_4_lut (.A(n28484), .B(n13621), .C(n2897_adj_2189[24]), 
         .D(n38222), .Z(n2937_adj_2113)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam div_13_i1923_3_lut_4_lut.init = 16'hf1e0;
    CCU2C div_13_add_1847_17 (.A0(n13624), .B0(n28462), .C0(n2699[23]), 
          .D0(n2641), .A1(n13624), .B1(n28462), .C1(n2699[24]), .D1(n2640), 
          .CIN(n30980), .COUT(n30981), .S0(n2798[23]), .S1(n2798[24]));   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_add_1847_17.INIT0 = 16'h0e1f;
    defparam div_13_add_1847_17.INIT1 = 16'h0e1f;
    defparam div_13_add_1847_17.INJECT1_0 = "NO";
    defparam div_13_add_1847_17.INJECT1_1 = "NO";
    PFUMX i32500 (.BLUT(n38407), .ALUT(n38408), .C0(n63_adj_3), .Z(n1351));
    LUT4 div_13_i1112_3_lut_4_lut (.A(n28562), .B(n13640), .C(n1709_adj_2169[31]), 
         .D(n1643), .Z(n1742_adj_1423)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/guilherme blanco/desktop/college/embarcatechfase2/placafpga/projetos/projetolaser/pwm_led.v(75[19:46])
    defparam div_13_i1112_3_lut_4_lut.init = 16'hf1e0;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

